��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�\�� ���K�O�{���b���ND��>N�!Kc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<�w�>��S�Ś��
��H,7!!?�#�1�:�Ω��{:R;ޒ1 T�V	�tL��	ǖ|�NiUR!�`�(i3�q�9�ͭqt2�*�����-�/Q!�`�(i3!�`�(i3�1B��ӿ"#~j[O\�K�y؄@�!�`�(i3i��ԇl2�����Vc�r5�:�!\Vn�w;J��w�4
>2�����Vc2�����VcJ�g�Hغ!�`�(i3ؤ�$!Ѫ���]6'�u2�����Vc2�����VcS� ��y�t��|���2�����Vc!��.���j~����B��S3��V1֛s�ӱj���fI�i3�������8�e$�1�D���")�/K�L���\��2 ���J��&�S]���}��U��=�A�PvH���mwWA���c�0�9���K��S���9�Ec��H�>)67F��UH&��p�M��Z̸*�����&�SV��"����R�i�cC��D^W��|��0����WE��/���h��p�f"���r������4� _;��i�1],Aبs��0�}bک��?���)t��⫓���3B�Hj7�lu~�~�y�Ap�1�G�$U��Y��U�W�8=�V����8ɞ�mQ�Tr�>b�L]���}���h?���+�t���P�����-ӅC8J���_NUl��FC�쌓���ew2�\��M!�nz��m��+@ˏ^ow�Y�`�o`d�kN���9�ĒTC��0���M�<lbts�I�Λyi�ZN�x�w�>��SU��Pa���PPe7m��������n|s�)>E1&7W�$J�|(�����	x]�<��O~��������@���0f�*C�"�L��v��d���.���X�����]��#���X
� �AH�ah5J�M��
��m6g��A� �oQx?F#��_L\�Յ�B�֪��Gu���h}j����5T%p5U\�����	x]̅���OI�}c�J�M=�-ě��G�$�5�	�s+џ�_�v%�L��xE*?V����
� �AH���CdZ�G�u� �(��Z�N��\�T�ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P��\�4�s��u�@�
�ԟ�d[u����lf/����Sd,�ϱ�)ů*W.Ӻ�bl�k�]vX��J���{�Z�JQm�!=�y����h�}�)���32ę8�����8-���/���Sd,�ϱ�p�`����j���$5�?� �٠FN�[\�i�]|������)*�M�����V�^�&�����!ښ�m��<v���ٌʪY�����iUM?a9-�7-ڍ�qL�\�X���щ;�a�g&C�V8����0�P.!܃��L~΄gO�3�:M7bR�u��w)�S�5� �7��Mv�9*���f��^.Ğ�	џ�_�v%�>+�$�~G�6֜S��0 ��D�W��.~�٭�Jر�D�8�>+
� �AH�)��H�� �b5z��j1�&G��	�����ロ�*�T������|�OA�
܊��?Y2���3")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F��_���P8Ad��q�G�+��T���jB�Fg�Y씤`��p}RQaI+k�U��OV@������,��B	hI�ˋ���'M��j�*ʹR.���U� ���_�o�ǲ=G}���@/�k�w��-zL͊�q��� ���iQ�J�x��|Dr�$׶��b9����4�6�t�����\{8����\.Wl0��F��jT�����N��>`�8�ux�k�-6G~���M�h�k7=����)�)�qT;l����o)�]r��*�S#�b9����s�AJL��<�!�d�<���9�����?�!�`�(i3�����5	���]���>����C�Gظ0����!�`�(i3c��Et��q���U��>�w�Y�#���\��Fw��|g�Y�'���Xw�j�7����w�K��ݑ�][H5���8�R�wX���c#Xe�l�`�B7d�N�By3��<�]�!����M[��ǢÕ�=��"�,�>E����-��%Mό���.�A�۠���AS�N�By3��<�]�!����M[��Ǣ���+1��;Ai�Ő��-��%Mό���.��D�����.g"}�p��Yl���#�]�!����M[��Ǣ�K�&�a�Ɇ�������-��%Mό���.�;�~��-�fu.$���N�By3��<�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳����^��φ��<�6�#b|���Mc��Et��q���U��>�w�Y�#��[H��p�����5	���]���c�A�L' ��a���R�wX��>�Q�c6���[H��pYl���#�]�!��	Ǹ�y85�����3�|#9���[�	������Cs�]2�y�Z鎬����[�Rs&�gg�C@,�d��E����F7G#+��\w��0]���q�D��`�B7dԘ]2�y�Z鎬����[�Rs&�ggλe�9�Č�E����F7G#+�Ǘ0z�cULjaGkƊ~8����\.W^�V]��}R�wX�շ9lD��XHӅ� T���Yl���#�]�!��	Ǹ�y85�B���0�1���U�<�o���8���/��,bxqX�z��W�����.}եӹ���ã0y���R��Eq(���#��C*�}Q�'����Y'��@UC��M���'�<��a�X�c�S��bƬ����
L'���Xw��e��c<m�
���n?~Ll���@IE�U��>��l%i�-;�ƽ�/��e޸XhZ�����
L'���Xw�j�7���S�ڬ��M���q�tt�g��U-�eaԗ5��C��U��_D��.V&��B֥/~.)��3\�R�F*}�c}��uO�Go@3w�^������h��Owq�Y&���#�{�0;�}����\�w�Y��k��ı����V���}���s+���#�x���c=��P�x��r��VYW\�'g`$�Y1#��Z�����XP�����w�K��ݑ�][H���\Q^���0a=cj<���|0���)ÒPl����u2�;Z�g��z��%�/[����n�[I���i3�|)sՀr,��>T��M��cg�P�z ��y�����,D��c2�'v�]��T�%q���IMdK�Ch���d;������Ga��H>+�w��0z�cULjaGkƊ~8����\.W^�V]��}R�wX��}�
�?�X����_�2^��R#��]�!����w�Հ�z���Q�����8��T��s�N��ό���.�c5�e�%������6P��q����R+w�7�CBg�Xs=��n`5�fK�\w��0]b!��u�=7�7K�P���������q���U��@����gGXWg�CTg�z�&��Z鎬������_�,��LE-L [�W��L
��JHn��z��ч��,1��; |�$:�c���s6��ݓ��E��*ZV)�J3'T��߷�d�٣��c�A�L'ϸ��%\A�����?,0=]^	�&|#9���b!��u�;s�e�$X�I�K�9f�7s�9���o>��l%i�-ݓ��E�e���F�&5����'���Xw�j�7����w�K��ݑ�][H5���8�R�wX��}�
�?��T1�8K���A�D��n`5�fK���ġC��׸@����gG�6�!
����"����]�!��	Ǹ�y85�B���0�1���U�<�o���8���/����,Dʝ�o���V��#��6��Q]� _ό���.�}�
�?��`�mp8V��%�TgR'7s�9���o��S8�<�)��'��*�S#^�V]��}R�wX��}�
�?���m15sV��#��67s�9���o�jƓ�[b!��u�����Yj<� �1��d�٣��c�A�L'ϸ��%\A�����?,0=]^	�&|#9���b!��uፘ��|�~��F�Ib��)'���Xw�j�7����w�K��ݑ�][H5���8�R�wX��}�
�?��vW(�������<7u7s�9���o�jƓ�[M�|a)� ����35}jQ����4|�����b��!�qg>1�Pq�@\w��0]b!��u፽��3rn�rMVXP�'���XwI����"�;�7���c�?��Ϭ��'���Xwx�����(�F�ܓH�;G+�ه�ݮ{�30�����ʍ��зq8�Ј'���Xw���,D�
�eM�6��`�B7d��n`5�fK�\w��0]b!��u�7�UyR�j�=l���]�!��	Ǹ�y85�����3�|#9���b!��u�s�Uo������zL�O�]�!����w�Հ��I��JnSl{�]&"(���+�J���q���U��@����gG5m�E��P�|�Ȝ��7s�9���o>��l%i�-��s=q�SbK����D�7���`Z鎬������_�,�����?�!�`�(i3%Ah�%4
>*"v%)��2��������� +_�XF�%�/kѶ���� ��Y�����E����F�'n�^0o**�ХM
�nGZ��JP��8\�S�.}�
�?�Y*�Ld�=�������d�٣���N N�S�qg2�K?\|iQP@�I	зq8�Ј'���Xw���,D���S�!�`�(i3�n`5�fK���Qi��+�`�������H���,>$�p�{�㘽2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��$O�a��Q�ڃ�)oY��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcZ��O��<�"��~Ǣ�)�s�ި�/$�ߺ��]�P���Qi����$~@퍜��Y�ؼQn!���Cs�9�+��N�5)��Z^S�QQ5��:ux����7��f:���x��
���Va�%��jq��/�a?�Ҟ��wɟs��A��e�����m�(1���&�����wɟs��Y�b�ν�r�� ��*ZV)�J�z0=�_���T1�8K��}!�#�b�Zj�|���ghR�P¢	�B�d�ZtgQ�9OZ��Q>ml�,"�x|ٲ��I����~u�g
�t����Zj�|���:�rQRт¢	�B�d����ψ/�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-�����*��=@rTnG��Q���;�Ӏ����QS��N��̉���G�+J��d�,1�!� ���үA,�&c����Q�nT ��{g�z�È�/&����� B�&"3݇F1�k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������7�,��n6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G7�wtMMP�~�9!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�Y������-JF����c����F��O�\E�W��4b-Ukc��R*SƇ���P_�2î��
�Ƈx ~����Z|
�Xy|�W�8�QeQ���{�`b+���Ã�-읟����u�H�h-) �w� �� :b/�Ti �P���R�!�`�(i3�q�9�ͭ���D��U�����i?�z�&Q�TyǨ�L:�싿�<��k�� L|��(�!�`�(i3!�`�(i3�7uw��8�#4�?�G�{�`���φ��<�6�=�Y��q�$%��W����' �Ϟ)��K������f9�&U�)j�S���ܚ��@��f�\%`>��s�;�jmT�#�0M�Ŷ�Eʨ�`N/������&G!�`�(i3D'm�����Z<��A!��,:&Ȍ�g�F��6x��w����Q�TyǨ��A:N� ,IİB���_�٪�(BZNp!�`�(i3�FW�DVx>74/���S�%�[!�`�(i3��b��~� :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3�;Si(�����_j��� t��RYr��}Dq�f��	��x��ݚ�Н�jCH�d*��=����h���ʘ׋�\!�`�(i3���F��O��ݚ�Н�T+���f�ԬQ���Kͽ<\��1tSjv�9��n�7�Y���_j�����9�x�\M�ݚ�Н����F��O�VA�ڦ�c4�f���^�
�3��Y$�VZ�ڋ���Y��c+�b�S�i�H�������+1�;�.��1���-����!�`�(i3�ґ`�g�y z�P���[���}��M�?L}�7�n��<f��5p�T�ۮM���y��C�o��vr5�Dѯ���-����!�`�(i3�FW�DVx>74/���S�%�[՝� s�#t��ۻz�˾ �����]M?��y�!�`�(i3���ܚ��@��f�\%a�ۊ�0,B!�`�(i3��:e �>���F*8k��.ͥ�H�RtV�^CH$�I��*�M/*�3�F�N��9R!�`�(i3��Ě�����}Dq�f��k��^�1���+1��*Hx�g���-����!�`�(i3Y�5�n����N6�������&G!�`�(i3VZ�ڋ���Y���GiL�~�
�:qEp�gdq�_x�ֺq٫[_�mS8<�n�ݚ�Н�jCH�d*��=����h�TGaG��7�!�`�(i3���F��O��ݚ�Н����F��O�VA�ڦ�c4:�!��P��3��Y$�VZ�ڋ���Y��<�{����H�������+1�;�.��1���-����!�`�(i3�ґ`�g�y z�P���[���}��M�?L}�7�n��<f��5p�T�ۮM���y��C�o��vr5�Dѯ���-����!�`�(i3�FW�DVx>74/���S�%�[՝� s�#t��ۻz�˾ �����]M?��y�!�`�(i3��#�a�Ąp*�з=a��o���H�RtV�^!�`�(i38�����FJ74/����1?�B���!�`�(i3�FW�DVx>74/���S�%�[!�`�(i31���~!�`�(i3VZ�ڋ���Y��c+�b�S�i!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 ��̢k����0M�Ŷ斗���%�������&G!�`�(i36��J��c�� �����]M?��y�!�`�(i3���ܚ��@��f�\%�~��\��8!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��/�"����I����޲��>e�FW�DVx>74/����1?�B�����#�a�Ą�ԬQ����5��t�1tSjv�����l��Cd��9s��vr5�Dѯ���-����!�`�(i3�FW�DVx>74/��� �!O�Bl!�`�(i3��Id�!�`�(i3m�����G����-J� �J�l_�j����ʉ��%>�rGO�D mWN՝� s�#�=�U�u�íN=]8k��.ͥ�H�RtV�^pT/�GS�7s5kL�G��Hb� h�ҩ�9��n�7�Y���_j�����9�x�\M�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 �t�td���5���d#�����"k�jCH�d*��=����h��LAи�����l���KyX�X:�^ao�&�U��f�!�`�(i3}I�6���N�Cٺ��G��Hb� h�ҩΪ���l��Cd��9s��vr5�Dѯ���-����!�`�(i3���ܚ��@��f�\%`>��s�!�`�(i3�k��^�1lv0�9l�d9=���u��r��!�`�(i3�䉌�+BNp��['���ڹ	�md�'o0Q�N����6 fd�i��z�����$���n"l}΀-/߅!�`�(i3�|����� F���du��1V��9`�p�0�R�y�����̚������Q=�ݚ�Н�9��n�7�Y���_j���(��2`���ݚ�Н�fĉ>99��A0ok��
�:qEpj�E}4ظ�N�Cٺ��������� h�ҩβ��y��lDW�Ĕ�VY�h�^-�q��M�$ci���{2!�`�(i3��w�`L�ķ@���k>��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t`���*1(*�O�qe��0�U���>e�FW�DVx>74/����j�����`���*1AL(�z��?�t�ϗφ��<�6�=�Y��q�$��9�"�5�:
1���Ƴ��d�L��E�u�N�iK�D�b=T ��q�z���v��6Z���,�,&�eǦ�@���<��+�R�`E�p���%�T����
�I�E�eNzL�h"j�j�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3jj�An%��íN=]b~*��s�
�I�C��ށx֤�%�!t)�!�`�(i3���D4FF��&l�--|iQP@�I	��x���^�Q:��Tא �k/�ݚ�Н�!�`�(i3T ��(՛MSc����h��N�M�uz�M�Ӄ%�K��^/p#��I2�8��[�@����`����ݚ�Н�!�`�(i3�����zCݮ2�����(�O>�rgBOY�]y�a�����o�u�/�tL"[$��$���ş����c�d���=R�.���#�&˸�rk!,>h2&�\0=��d� WF������ɐ�c,h��ws�M m�o?��Uv�=����������Cݮ2�����^���u�s�d�p��<��wFB�b���t�T��?E-h��$^(?��"]�B���[�.��|ȃ�A(�c���_G��Hb� h�ҩ�pॻ}��$�2p[_��dN�<@Iv��nt=:��:5A��p����g�Z��3��a���!@�f")u��r��&�	o���,�,&�7v���Y���+1��*Hx�g��a+�߅� �����]�?��6�=7!�`�(i3@��	Ķ=�����#��[��o}��,Y^�{��b�b�*�����u��r��;�~��-�f����Ga�߈.m��B��+�T[nHN��R��bP�63Z�t�5ߧE4��Fr��j�:����|_e=���s;[�T�����Z���6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G���������'|F�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^[�5���78�íN=]b~*��s�/$�ߺ��]���޵.��g�d�H�RtV�^�,�s��(X��*H<s)l໶�,3��0����[��o}��MX�w����D�����,���-����!�`�(i3%w�*�7���?��۳lU����Ga�O`�� \)��w�w:�!�`�(i3;[�T����kb- m޺P��l_��H
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�^�#�nish�Ž�������"��T��Z|�M�,!hޖ�A$�P������5d��n4s1�U��B��-3��܌o�_/�2��<�7�癆cgQw�c4~Nr_�mS8<�nhDJ��3�~�+yp�l�#QSU:��8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�/�e�i!l��íN=]b~*��s��(R\֎u�Yd�E�WM�v�?i�:!�`�(i3&�|Ξ쭔|�~��ӂ�=�7�'��ڎC�?�x��w����֯���,mk��L���n��<f�`u0�F��a�7��]�ݚ�Н�U��p��PrΌ^pG2��$�)�vx�;�U4�Iȗ۰�=!�`�(i3��j���"&yf��o;��0~�$�q����ڒv�4�?zm�X�R&cE�����"ɻ���&@֍���,�,&�X��X%�B�`u0�F��at�zEw�7?dq��!�`�(i3���3rn<F�ڴd0��d����"��
��h�/�f��Qc��Gx�˔��� �So�M�{��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=��F,��C-[�M��Ra])n#���r����)�{6�U���[�	���d�~{��)P<�ܓ�Yfĉ>99��A0ok�����F��O�\E�W��4b�^�#�n�~�+yp�l@�ߋ��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��N��[r�&2��m��)��^u2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0l�x8��-V�s�u6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�27���^�R~T��æ'ž1�|�'����u��r��Ư�ճ�%6�E~�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^7�UyR�j���;��Qe��0�U+�qbp@�;�jmT�#`&c�'N�j�ڎC�?�M?��y�!�`�(i37�UyR�j����^7���!���e�p�x��;b�-�2�ݔ�(v3�l{�]&"(�'����u��r��>�Q�c6��=�ڹ&)�\��H���gY6!�K������B�̢k�����U�R^p���P#G��Hb� h�ҩ����q�D�-c[����K/x�]u�
@!˥�I:��q���Ě����>=:9_�a�;�P�t�5�׹�� �ѕC?",I�$�*�����sdJUX���˫φ��<�6�@a� ��fFMqlg{y����i�q,?5q�ӫn>�!�2G�,��R(bs��2[�a��o���H�RtV�^"��
%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���r5�I��d,ܓh�,������&G%?gV��UXi�G�y��״$(�>g�fĉ>99��A0ok�� ���Aؠe
�M����d��-��!g��J�s��z�
1���;#o�]�ʄǝ��pك �%�K��^/p#��I2�8��[�@���=aS�H��ݚ�Н��&��>��q9+t�}�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��&��>�@�ߋ���|�G��p���~Qy����?��~g���C>i���,.��uݑ�4>
'�=���ۉ��K�M�,!hޖ�A$�P������5d��n4s1�U��B��-���忔8��;	ȕ?�7�癆cgQw�c4~Nr_�mS8<�n���*y}e�߿�wW��C�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�`&c�'N�j��O|���/��kOT ���Aؠe
�M����d��-��!hr������c�����+A���:�Xu��r����Ϟ4�>Ht�u�Un��뾦����%>�rGO�D mWN��Ě���aT��3G�IX0F�Ms�Uo����N6-	��6<���{k�˖�x�󢯖^��'�ZT�����sz`F���.��n��܆���M�,!hޖ�A$�P������5d��n4s1�U��B��-���忔8l{�]&"(ShT���A(�c���_G��Hb� h�ҩ�`&c�'N�j���$�a/��kOT*qA����6\�4�@�� �-j�1tSjv�œ&|�9�n�o&uL�)P<�ܓ�Y�H�������+1�;�.��1��r5�I��db�W�
�a�	�Z���ވ��*I���b�Bϱ��>1J���� ��0� 1tSjv���(���0�l{�]&"('�^�����;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�`&c�'N�j�ĥ�A��o2Wv^᢯��0��鯣��PSMǓߥ�{�w�],���zn��!��h���ad�~E6c�s�9��᢯��0��.T�Vَφ��<�6�@a� ��fFMqlg{y����i�q,?5qxŴ�Đt�|�Ȝ��ShT���A(�c���_G��Hb� h�ҩ���U�R^p���P#%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<�a�}�$�᢯��0����$�a/��kOT ���Aؠe
�M����d��-��!�Ӈ�<�H z�P�����+A���V��𕛺"����0��e���F�&�?\MP!� u��r��w-)Sz�M�:�.�N������4Yz����|e"���F��O�}�	76�&�� Ӗ�t$�)�vxկz|h,�`(�w}�eX2����Ɔf���l�����t�T��?E-h��`f���sd�G}%����3f�m����2G�,��R(bs��2[�a��o���H�RtV�^��S�V� h�\��;�,*qA����6\�4�@�� �-j�1tSjv� ���Aؠe
�M����d��-��!g��J�s��z�
1���;G��Hb� h�ҩ��)��S�2���i�AԢ�a\�2}$#h6��8{4����gs)l໶�,����l����iﳇ��� +'ێ����� h�ҩ�'9�и��{����@z\��}Dq�f������!�`�(i35i�a�vb��}��;�b��~$�
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b��Q+��
ŧƧ@�Ezәߴ�)n�?M�,!hޖ�A$�P������5d��n4s1�U��B��-^;�Z�N��ShT���A(�c���_G��Hb� h�ҩ��j<��?��;c���k+Q�h'�Ȝx�5W ��̫(� h�ҩ�6��J��c�eK�	�$V�G��Hb� h�ҩ�|D
�W�ɪo��<�����	G0��t�UW���.6��"����u��r���"�чE4�]�p� �!�`�(i31���~�B�'��a��;��%���b��~$�
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b׏�����-�5k\u����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h/KuTШ�?��	`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc ���v�[��|�z�|���{�G�!��A$�P������5d�	�+�&I(&�L��'ž1�|�'����u��r��[J�2�����瑃�dN�<@Iv��nt=:��:5A��p�s]��z��(ǝ���q9+t�}�|#HK��e޸XhZ$�2p[_��dN�<@Iv��nt=:��:5A��p��m15sV��#��6�q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK���7�^t��d��-��!g��J�s����0�|섃Va�ir{��b�b�*G��Hb� h�ҩ����\��(ǝ����ч4H��&��;�t/����>�V��#��6ӄhD���� )�(��!�`�(i30: ��qx��c効j��
��e޸XhZ��}Dq�f�n�(&�)KYO�*�q ��]���
 v=}��a��;b�-�2��;�P�t�5$f��_Ub�,�"���M߸��S�Ȍٽt� $�N�]��V-[!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�x�\o@��L n�ݣ�`2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�w܊�r%�e���F�&M�,!hޖ�A$�P������5d��n4s1��7�癆cgQw�c4~Nr_�mS8<�n��=����te���F�&s��>H�,b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vNd�8��k�Ss��Zf���g�F��6�	�¥�S`/�dI{�b~*��s��J�'Ƕ.XC������x��y�o�!�`�(i3�>1J���J.���\f6�i�|?���߆�p�h�՟,�tpzuʖ3�z{φ��<�6��`䘸�|������&G�B�'��a�e���F�&G��Ye8{b	�fƏ���%>�rGO�D mWN��Ě���aT��3G�IX0F�M�>1J���W �8�j2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�h�V8�&FY0Ƭ���IT*O�.2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc,I���H��Y�b��P(#yc�Q�o��_�Rv�䩲$��8��I��.��|ȃ�A(�c���_G��Hb� h�ҩ��T1�8K���A�D�%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�m���>#o�]�ʄ�M��,����q���f�e�x��w����֯���,mk��L��q���3�tޙp���/�dI{�n�|�-3�A���|���d��-��!�"ǉ�t���S`5�㬌�$Q� �H�RtV�^;�ƽ�/����R#�K�|�g�.�n;c`3jYYf՝� s�#yM�j�PF;Ό^pG2��$�)�vx�;�U4�I�';��#j�ݚ�Н��T1�8K���A�D���ZY�ru>%L.�A,��}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ���������zN�S��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Y�����}Z�
d~� +�i;\E2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�p��Ik|�Tr�ҷn�^N�=���G�@���M�.� ���ѡ��}Z�
d~@�7Q�wm���7���6��&�(\� ���U��s��6B	�?0�m��I6�X�,4�?n�[$��Q�h��*
ak��h*-�#���~Qb͠�Ԏl�>�xj%�;'��V�j#�{D�A�W+��W��`��&0�yl�q�����U��)��~0&ۅN,3[{���:յ[+8�SݳD��zJe޸XhZE�g�������(ӈ���m�r������=�g�H�:��a=�9$[{^J����{J��3	�o�{��q��"o'���\�B�ݚ�Н�r��Ɉ�?����2���N���!�`�(i3����SP��'�K �_�mS8<�n�ݚ�Н��7��aM*:�b��t��������\A�����?����S��V�H���@��i߫�\K״$(�>g�!�`�(i3���F��O��ݚ�Н���jVѭ@!�`�(i3i}B2>�~ �<j�"�AM?��y�!�`�(i3㣅Dy�'0: ��q�ˬ�wO����b~�>H�U,V!�z0���6<h��?D�8�鉅�%>�rGO�D mWN���%>�rGO�D mWNHN��R��Gu�"�0��Fr��jj,;P�j�w�R���y>��yС�&�b�j%$�^^4>�D�j��A�0: ��q�9�|�k7 �@��աbR�I�/X�
@�i��g�?�d���&�V��o5]�:�b��t.�C��6�o8:4ښ�*jl���C>��ӚH�RtV�^����Y�z0=�_���{_8�Y��=�}�Vݨ��}Dq�f��R'cf��>��YfG��-}RY
xǍ�J�r��ps��u1,����Uh1�[��(��;�jmT�#PB��/���߰�$|�Pu��r��;�jmT�#��	�DůI�߷�c/��-����!�`�(i3Jº�FO"V'PS�����S�ڬ��M�kDu�H�f�#��(�D�"��ӌ�r!�`�(i3�5ߧE4��!�`�(i31���~����l��Ht5�=�5����������&G!�`�(i3SݳD��zJe޸XhZ��-����28��m)�+#��E�#Д¥���|e"fĉ>99��A0ok��fĉ>99��A0ok�º��W0�]��x@���׹��L<C%`����,�ǰ	M,��rER:�b��tu���oܢ]���#�;¸�[�E�ȹܹ���8��<G!����xQ�aY�ix�P�R���Jm�W<�WCۓj*0: ��q��+}�_�U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&GK��ft��;�cM���/.�,/j��O�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�ґ`�g�y z�P��	���QC�íN=]b~*��s�/$�ߺ��]���޵.��6��t�b�!�`�(i3A���|��`�Y���p�_5�?*���S`5��Z��kM�8�/�dI{�u�>Y�u��r��9lD��XH:�b��tv|	C�������Y,�֮�Ra])n#����!��:�8QG8�]߸��S�Ȍ:�^ao�&�U��f�!�`�(i3<���d1x��r-�T��y��BQ@2X��K���q��Ɨs$f��_Ub�F�S�1 �;�V&S�bO�D mWN��ܐ�}Ħ8��f�+0: ��q,�9��!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�v�����	��Xx����Q��T�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc-�u�b\�W�X��\M��T?�d9��AdF�����'i��'�I���5�T�U��'"!�U��)��~0&ۅN,�~ޥj�!W�.��|ȃ��"B��XY�4�A���Le��0�U+�qbp@�5�����}Y��	}�@�im�1:��am��	t?�*|�c��>X���4��G�)[7h���;�jmT�#PB��/����ƾ_�u��r��Jo���j� ��7P��'����u��r��t����}�vߝ��y�b$��o޷n��뾦�!�`�(i31���~����l��"B��XYQ;1�'�3��q9+t�}�ݚ�Н����F��O��;b�-�2��;�P�t�5���W0�]ݽJ/��v�$�)�vx~�O@�d八����T��_�Ι2QX�o53�_�3�����|�~��m�G�V���R�m!	�quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7�)��yB!�Y�(*5�Y\���F�`yx�>�+X�M?��y�P#+_]ݱ�x��
����#QSU:��8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�D'm�����Z<��A!�!*��*8�N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s��ݚ�Н����V[���*φ�\-�g�W��L
����LG��&{��b�b�*��7<M�u��r��9lD��XH�H�߳Mk� ���c��9��'���߆�p�h�՟,�tpzuʖ3�z{φ��<�6��`䘸�|������&G�B�'��a����w���VŬ� ҿ����qJtW���b�0���Ě����E�i�m}6O�D mWN��ܐ�}�>]6�����l��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc҃ڹ���@�*�>U|'2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�j��A�<Y������q8h�9MHH�7� a⣃_BR���Bk�dQ�TyǨ�%u�X%��d�bB����\��q9+t�}�d�b��6�a��)P<�ܓ�Yw�R���y>��yСs$8��ѡ�X��B���Fkbҝ��q8h�9MHH�7ḩ��H�V���羹��`c�N���GedTlya �x�x������w	}��SڣE�,E9�1f��P���P,�ǯ3�4����%!-�;������ �5p�T���w$�tJ�rS�b�8Z�AԢ�a\�2}$#h6�� �4�u��XW�����_qa��P�F�|���#�ҵL��z�*�&ƃ��#���+.f#�\���Pi�-��M]�5��U_��{��b�b�*��x���_nY<�m��Z<��A!�!*��*8�N�Cٺ��#o�]�ʄ�߸��S�Ȍ:�^ao��
n�Ț�)��b�Bϱ��LU=����QY#��I2�8��[�@��OߙYĸ-q�A��Д1���~!�`�(i3?Q�@X>#�Ԥ�8!7=$o��ɝ1M�,!hޖ�A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�7�wtMM��6�a��)P<�ܓ�Y�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н��� �.7�|ʓ����kb��H��n�-:��;?��Dƺ �X�[g8@�ҭ۔�P��V�N�,�}��	�8�T���y��lD�6�B7�� �3���=�B9ٷF�����l��$&��(��t�;!��QxP+�L��k��������d9=���u��r���#�-�p�G�6�!~�%��v��!�`�(i3��Rx��ڎC�?�x��w�����ԬQ����5��t�d�8��k�S���ȧ]���b�Bϱ��LU=����QY#��I2�8��[�@��OߙYĸ-��-� 4�+D���Q؃�L�\�@����_%}i��w�&�2���������!�`�(i3	�%��6�X��ͷ(�-���|e"$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��4�5�$S����N�w�R���y>��yС �ݻ)�9µE��\6�5d�[�IX0F�MV�ҁGG%4vkz����`���φ��<�6�B䁒_[�FShT���A(�c���_G��Hb� h�ҩ�B䁒_[�F�q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK��$&��(��y�`��vN	���QC�íN=]b~*��s�/$�ߺ��]���޵.��_�mS8<�n�ݚ�Н�B䁒_[�F'�^�����;b�-�2��;�P�t�5�H����{��b�b�*������� h�ҩ΃�f�,�k]�(�����!���|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�?.8h�.�z��Iq��R���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�̣n;��6����gɄ�6�o8:4�I���c�90��G��6�iI9�o«IX0F�M
z���\���F�`yx�>�+X�M?��y��#�-�p�W$q(W����?D�8������g�Z��3��a���!@�f")u��r��%�r�����5)��Z^�'����u��r��N
�����"ª�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��N��)��V�N�w�T� �f&���#��D<V�-�b�+�