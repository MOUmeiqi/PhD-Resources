��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag����pH��q�P��'�<7\F���r����&$9g8�M>PFWD#�z":���ӳ��_�x�$t�`a\�R�F*}Ø���K�ZF��W��`k�ZV"���:��#tC���,?a��Q\�_qť��[�޿J�F-p�-� ��d�n}K-J��K��z������3�z�ω�C�I���7��@��	F72��{L�8br�.�/�d�������4�;���u�$|�>I��4�Y�YrT�#.�Ő�|��h����jǎX������n�q���xP��t䗒�|'r�tI����j�6ˊA뫕p)1 T�V	�tL��	�<�A�}Q@���rahH.�J#B&ljW�n���8�U��]>��D�,�Hc�.[K��m�X�'b�mh�@� �ʁ��+��| '���贅�����OW��F!���p86_���Ӎئ��f%%e��h&9�4[f6<%L����d�؏	�U��Mm�)|O���3�dR-��S�0I$�o�W{��ǖNfDKA�1��xL������s�3NX������1Q��?�4�ʗK� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F~�?|�[_wȵ�e�kY��Y+]��tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Q�{���_��Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��P��'�<�磋��w.V&��B֥/~.)��3\�R�F*}�c}��uO�b�^��\/ɭ��:�Rh�&�~��ea�;y� ����t��!k@���v~��<
DN�!�`�(i3�b9����$�n������B�K�9gP�U,��!:��Ok��@zL͊�q���]p�Rrp2��ͧ�p9+�8��)(j�9v)�Dj_Q���V�Ɠ[v�Bx!�����m������
����:߀�����9��A�����y������i�!�`�(i3���D	��U�l>o��|�,+$\�M�ƕ�mo�0�VC ��0|]<w:�!�`�(i37�ܥ��2����*��5�V��On�/����Ʋj[�YP����M�g����!�`�(i3�E����F��j��\w��0]瑲��Zr�zM#��m�"�,�>E����-��%M�:2QYeƈ״$(�>g���0�&�ͭ�h�O�0"�,�>E����-��%Mό���.ӏwbk�$���7Z��!�`�(i3c��Et��q���U���
��I�PM�'�ghR�P��|g�Y�'���Xwd�n]N�/��A����Q[R�7J���hB;��i|�l5R�E����F��j��\w��0](@X~�H:6����Z9"�,�>E����-��%Mό���.ӈ�=�$��zigzA=v)!�`�(i3c��Et��q���U�ЂDa��(%װ$��_�zM#��m������
L'���Xw�P���w��:
1����s�!`��z�]2�y�Z鎬�����	�7 �# �����2�w�����|�Ƹ��]�!��	Ǹ�y85�����F�>R�wX�Ձ��̰�!w���B}s�!`��z��(�
t�ژq���U��d�b�ʪ%��1!�`�(i3�����
L'���Xw�4��}�<܊�,��!iJ!�`�(i3v�ј�"��Z鎬�������(������ҹ����lC��U�T�\ ���A����'Vp��U�!�`�(i3Yl���#�]�!��	Ǹ�y85���~iI�D;�¬pX��g��U-�e�,���6+���&��Ө�i|�l5R�"B��$I��w��,�񁫴}2��8X���4bS�N1�	(f�`��2&+��T���jB�Fg�Y씤`��p��>�B��7���
��D�#�U,M� ?ҡ���y�E�nwE��S��q�P ڨ���"kA��8Z�ZVq+��T���jB�Fg�Y씤`��p��>�B��7���
��D�#�USy���5�e`��9�����kO!�`�(i3��Q]� _ό���.� ��h���uT	���!�`�(i3"�,�>E���]�!����w�Հ����b����U���g�7s�9���o>��l%i�-5�e`��9PB����AP�p^��g���cό���.�}�
�?��(R\֎u�D��u�(nȯ�?
YT'���Xw���,D}p$_~R�(�[�*"�,�>E���]�!����w�Հ�*��9W��8�����JC�� W7s�9���o>��l%i�-�u��Y'Gish�Ž�� 4ȶ>~!v��Q]� _ό���.�}�
�?�V�=���_���&#ݟзq8�Ј'���XwI�&�\�+1���}x*ؐӘ��b����/�:�3�TF
%$�����!���d!�O��1��2�.w[�%�!�`�(i3�i3<�f�D.`�Z���L5ӥ���98�
x�?�����tz|���~{�kѶ���� ��6@�$b0���]<���Ws�N"T8�zn6�u���Q0�lC��ۺ_~5�Ǫ��I�&�\�+1���}xe�4޸5b��F�)�}�����T��.��W����"�,�>E��ۦ� ~�p���F�)�}�����T��.��W�������E���b!��u�PQ�>\Ճ�I��b-���q�[���QR�hǬ�&Q���5r������.U��6�� �)�s�ި�p�m~|�օ�)�X[��A��:o384];ˍH���6��g�Q�q>x��U����N�b^X�P�w��9+���Y��J�y��*?(1#��Z�����XP���[|��;�W�x+Q�*a���]�@����gG7�6>ᙇ��5ǗcV�j7s�9���o>��l%i�-He�-�c��R:k�ڛ���Ο]_Z鎬������_�,��i�p��+���*��^.I��Q]� _ό���.�}�
�?����4)c-�¾L���d�٣���N N�S��E ����*{��[�$�зq8�Ј'���Xw���,DFmғO�4}�G���n`5�fK�\w��0]b!��u�<�`A��_i3i 
�c��]�!����w�Հ��a�e56<�!�9Az]\���+�J��Y�{'%s�:�f~=g(���B��������z(x��g��U-�e,%�0g��ա�a�e56<��f��E���$ r@{�q���U�pzl��a���8�%�b�-�#G�H>+�w�\w��0]��4�ό��r&����y{N�En�J�a$�Y ��Z�/�N"O��Z|)~��\������T���
!O:0����-yMc|`���k�����=ZXRY�bt�atbK��:z6j���H�Du�%ϔ�}��ycĢ���Υ�d[gJ�a$�Y p�YD<=���aR��E�K�&�a��aR��E%w�*�7�����'�}j�c�q�����0��G��e���������6~�^�[@�e���!
��D��u�(n���q���sv3����\C|0�����?{�������l���3E��ާ�����ݚ�Н�!�`�(i3!�`�(i3 [ad��ؤ���@����!�qg�XJc���!��{*9����*��� �iK�D�b=����LB�g�RMm�o���xӯ`�ح���i[)��V����>w�0�S�n�(�a���3E��ާ�����ݚ�Н�!�`�(i3�y��j��k�BT	��.���i|�l5R׾ŞWsuzPB����A���'飥�ƷD��kȻ{Zٜ=bf�й@�X�/^/���'�i�o�q�XU�iK�D�b=Uq,lLBP���aڽ�����C�#�,�IX0F�MV�ҁGG�K�BN
\���$�Qu�2[Y:,c��W��L
���d�٣��c�A�L'�����--��wء}��9�sN��ڂ�ޕГ����і\|{���0��iU[@� +�Z��~�vϸ5Eb�S;A{���f�%�2iI9�o«IX0F�M�ȏ֦�"�\���F�`y������T�8k��.ͥ�H�RtV�^%w�*�7��.��Ã�����ic)�̩ƍ2���l�J���hB;PB����A����;q��b+}y[�i+�ȕW��L
��!�`�(i3�ˇ�h��<�W�.�P�	��
�Q�}�%t̓�@�O����&{�A���Je��b+}y[�i+��_1�f���!�`�(i3%��v����l�^!�K�g;�UA�qIp��K����c
=^Lma��Ck+Q�h'�Ȝx�5W ��̫(� h�ҩ��W�3�-[)��V����I����~u%w�*�7�����'+�dr�����o�t��D��u�(n�D5���.p�YD<=���+���q���i+�ȕW��L
��!�`�(i3?����������	J�Q�TyǨ�W���>Ca(􆿳��3��TY�l�rx��E�x��7�֕iK�D�b=��p�:�S1�ӿ�Q�ЙMǿI?����[jMQ���0���g�����;q	�%��6�W���b�0��%t̓�@�8��"�7ό.R��x��� ��2�w����:��q��5ߧE4��i+����ak$5��f%%e]
���7������	J�Q�TyǨ};4lW5�CaT��3G�IX0F�M,yO�a�jmy�e��v���bQ�*�8������l��M���Jg]�B���W8�8J�|9155V�V[x!��G-�Xy|�W87�_���4)c�ݘ<�̆xڥ����Ⱦ��0�|섃Va�irD��u�(n���q���sf��V��y4k���Z!���Q�_��VF�˷��h��N�M܍�?{�������l���3E��ާ���虾�b+}y[ٚ�	.؉6T���QL����f����������֢&@��&2W�+�?"J�L�Y\ٿ�6�PC��uB&ǣ©��*��^�"~H�𕎭own�~]�g����A��`-�*������Э~���V��2
L.�X;p`��vbëdPJ�9�Q6f�?ǉ�=��R~�e��ד*�h��F�v�C�5�9�(��Vh��W��w�x�P���E�`JcU!�`�(i3XO����0¤լq��/&M���<�q��9wS7��_�_��Kp�h�x0�7l]�) !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��B��d(��.�����gRI/!�`�(i3�Y�M����4Wt#���MK�L̈́�vw�aS�>
!�`�(i3�M����v�v��8<e
.�Ūz�/>�"�Ax!�`�(i3��3�N;C�]�'X:��+�i�	��_�V!�`�(i3-��!k@���v~,��L���r�����bС
��!�`�(i3�X;p`���w�K���&v�`�L�eyk1hDJ��3	�_:iO�A��*/�|��&8�,�H*W��u�a�8�c-~���D�c�J�.��8z�f�h�\ƙkH*W��u�a�8�c-~��ԁ���T!�`�(i3�&8�,����0u�CM�&�mU�w�������*����	�?h���5�e S]#��+qѭ�+g[��MQNv�2!�`�(i3t�%�Z?�k���ҩrɗ{�� ��Y����
� �!�`�(i3��X)�:����s'-��hy��jX�p!C+Tl�������l6���퇇М1-�����'�u�f�?ǉ�=)�{� �"�X;p`��L�t��nf�?ǉ�=~n���,a�X;p`��B�+2�A�:JϮ|�秽m�&8�,��Om�"���^��Ɏ�#���?\a��4�czZ��������[�D���~�ߗE�%�� �-��v�-���w:7�sq֜�H��s8��!�`�(i3�$�~c/~�O������*������R���e�D�
�~��\��f��E��Ⱦʤ ����i�\!�`�(i3�$�~c/v��&EA){c)k�3�� ��L��4��Q�j�