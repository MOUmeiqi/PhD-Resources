��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR���b�z�>}��������q6N<��;���Z��4d��{�
��|��Ȋ)zo1���á�rezxB���]Zb@�q�*�+
MہW��K�F��1�:�Ω�[@�qR���b�z�>}��������q6N<��;��� B]�pE���	x]̃Dj#^Da����M�׍�ё�6ٕL\S��A�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��QՊ(�
�d?t���raУ�Ν��u����l�|���j8��6�ܬl!����Y�f��a�Z��V�H9�~r�}��%%��*��!?9(�S�E���XP�� +@�������	��c�U[�� Oag��Y/�]��ݨN��ggL�|�A]��3@Z�i�D��� i���u~V����v��6
R[>�y��W�y��MqZb��9���'7���	/ܘ���?�־�+��+ER���r� �C�-B��<���2O��'HY-��Yk"1/��n5R�%�.��.f\y㔪�_;2a��k���9�ĒTC��0��#3s�}�!#m^s?�������AEP�� �b U�X��o�K��>���:E����҇1���%[C	��}	�/yϻ�b޾wbC3���!��4�nξ��k?�N2)WasS�z�r�o�u�/��h_��E��W�0��q���Z�N^��"�ٴ��1H0}M,b�Xgg���[�hѾ��/@��<bg�'7��k�8���҆�|n����B�~O��YB��x-Y�lP���U�)�(27�׳�_�";Q �Ar���5�Y�w��'�i�xiq���Z�N05�����u��w)�S �J���vy��0ӵ4�ys���V�gL��˓f�+������R��j�EB�1~�����Ǔ?B&�� �=c��h˗�)!w�G37)�t��z�k���r� ʍ0�v��-R�n�Ar���R�G�)q�j��U�T(r�J�F���5GR?:2��At:�)6�+�!d���w
�`�!~�?�����Wu��w)�S �J���vy��@��."�^�S��J�^�M��v<f�+���:�8��?������
�r-����\ �?�����9��hMx۞�D��"�Y�
� �AH�B�5����Z�<uo����z
�X@���!L�����v���m)D:�l&����� ��t����dv��(�JR&��a��N�!V2T@\~�.���-���>�o�$��9<w�<��o,����]Iv4�YJ��qq������-���=a癪�N�v�ͥ�����u��w)�SU��T�d��6��.7<k��h��9/M�C/f�+���C����
4��YN
��)eZhpH�R�l��5�9���/A$TG�	8����J?1��r�O��C��0�����U����X(�7(�C�B��}�@�����]���_����J�UVN�����tf]ƒ��c�#ϱ����~7fx��zG܍�+�ł� c��(�U����	x]̸�A(=1/���ئ^��w��L���M�S�O1����E�`\��f��@9�¼�l9���ݽ����.��Z�������� ͗����:���c��$�-Y#дS��E%��൭��n�ZQ#�+��3p���u\����8��I/�6�}
�V[�W	�8�q> �:4�eȹY�����!ߥ�A�.��q�©������5X�/x��-w}�~������ۥ�A����DK�$s�B�+�V�p���������RL�a)�5DK��}��~篟|�<d�-n�L�FI��l9����E�E����}�c��_�+-�S�A���T�*�QKK�L5e������}0x��1�g~d��Z>b��m�!=�y����h�}��3��5kX�Z���k�W׉�oB;sѱE�DK�\�h����BPMF�I�	��U�!l){��&tV�O�����K����J��\�4�s*�*Vu]�Z�o/5�\ݶ�����N� �ֹY���8���+��"B`���^��G��OJ�O܏�M�C�D�~�&�o�i�$�NV��ݻ��3';~b����]?��R6Cm�!=�y����h�}��1��qFM=���u�2Ϳ�؍��oB;sѱEϪ��nȸSB�r��Ow���R��������]��)�HE�fśp�k�8���҆�|n�����ɬ��
�O_Q��fvЪ�M"���U�)�ΗT�0�!�g埿�G�(����i �ང5�}��S��&󑰑 �5��u��w)�SU��T�d���@��."���*(��m��X�BSf�+���]h�$�0d\F���+���\~K�f�R��v���"�9 \r�O��C��0��+J����:f4�������j���������\V��t�ee�}�]��]#S-3>��6~7_(y�,y��=�-ǺJ��O�~���RL�a)3��H���~篟|�M��4%a�U���y9����E��Jз&�6�f0� ���2�#�l��\�4�s��5��"�K+8�MK������b`'�$�ֹY���8���l[��4��L�5Z��%��@tOIkV�g��f%_�C�ʂ"�2��k�8���҆�|n���>������Z޶9��s�;U=)��U�)�hѳ�W�Ff�a4>t��ɘ<�-��@C��\�4�s�]o۬��K+8�MR�����蜓:�
LֹY���8v�J��f?C|�6|����J%�hu�՗Xr��ӹw�u��9�������R��Tx�&���jr�>,��� 5T��Ɏ���������	x]��r�Rby^K��l�Z�a��w4h��.*2SwS�O1����Vc�L}��Q ��<Ni�*�H��F�1՘y'��BS"�9 \D�GB<x��,�5��S��������,q�` v�%@ܣ����wbc����\�4�s��Иk@D��K+8�Mb����>���B9��ֹY���8�B�l��3 �gS�Ȋ�څ��h�7��sB��� e�P4��
� �AH�bs^&�m����0ӵ��Dc�)� ��`	�%îf�+���a�|goS3�M�D�I�;u��w)�S��X3�����Շ_ Q �4�=�z�Ǔ����~lf�+���@yc�s|+E��.5�����O�~N�G�}Ř&��E����8�
� �AH��%�i�6�K�(�Y���m�W cҝNߓ�G��L�����
��|ſ��f����1X(ݷ�u�0��bE@N��<b�jT�.����j���.�U	EX͇�,А�r�}���hv�(��z�j*��y����0��H��k.�n&k]���E�7/ � l�\�n!3�����(�^�K c��(�U����	x]�V�����K��l�%�G�;r����"m |S�O1���l&�ǿ�_\SEх
p+L�Mm�b����k!�\Z��K�������QѾ��/@��8�>r&���R�}vJ^�k��76���Y�Ɂ4
� �AH����e�1J����
���س(�0��&���S�O1��J�����l��Qr�ۯ�2�/�*Ư L�jy�����N\���&%�/�)��Ɍ�*����m��9��̵�%(u9��U퐑[�_�A��1k�J�`�k��?��k]m��C/S�*s��A �sb��E��@m�!=�y����h�}4�1[k�8�ɵ��aE#�����4���U�)�(27�׳�o+'�E}w���`�W�V��<��,��ƂYx3g�h�e}8�D3?@���\�4�smg�:�TZz�(�Y���m�A���$E�U�>��tL�����Y�F���)���@v�({����w"�W������RL�a)�G{�<���K+8�MN,�L���l�%�0���ֹY���8�d�5�r�O��C��0��`�R&.1� �Z��[H���1�<'"doB;sѱE�%2�}���3$�" ����f����m�!=�y����h�}��<]~8+|�Hў��͝AY�̉��U�)��T�e�8�޷����	[��ϼ���j�r�
� �AH�)��H�>,�
w�?��3u���&�r�ր�S�O1���9
��O�:�_e�"g�VƊ���XZ�D=,Ϩ4�R؂+�#感��{]9]Q]F��
2�h���'Q�����B�΀FQF�g"�u�̤�'�dX�Qo�n<�![0T&�F�=���Y�)��BĊ�K����*k�u��w)�SU��T�d��~篟|������JG�}���x�9����E������f�P��u�mw1m�!=�y����h�}�BK9�H�n�B�A[��������U�)�\8�4L�h~��(9��Q����q���7����3B�E���G� ���,_�kh;��FJJ��s���CLpZ�� �"�9 \:�ͮ�g��/8f��Jr�1��J�ahn��F�~�s�j�n����?�UѦ��	}����ó����.���5�y��z�qt4$p�o��'�Á�������50ck��W@�S6?���uS�@2m�ݸ2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q(8H�Yy٥;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"�"�A�-��ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+�/����E�{b�2"���Bpш�#w��q�©���B���������'Sea�8���`<4}��(����5��4�l��S5H�j.F��_���P8A��3g�ݜ��q�©�����Lu�m��+��$|��;D���J7"�"�A�-�#�̔"v�lf)@̲#;���(�s�-���f�i\􁗊�n��\v;V[���b�/ri�y�!�3]o��in�m��+�ڔ�wV���C�Sy6ג��̹��/R#�x���c=Ct�z&���t���Zu�2���8���Z�T�%$�����j��u��d��kq�1�U��^�ͪ�o��O��j���3�n�����j�0�B8�9���X�G��YG�g�b�+�y����o����+� ±�sR�{F;�f��X��a���x�yB�+�V�p�E��٬���M��҇+:|8X����\�v�r_���t�td���5ct�:��RE��Ok��@zL͊�q���Vǃ�����������-N���\�vņ�Q�]�ޝ��(��U��֜��3�b9���с�'sIP���1>y���Mw���1�Z���=���u*K6HT�����N ��S�����B7�B����{�����N�I4��欱���j���Ln��S�W�q	k���Agf�m�6��Rf�yoY�����-�h��7=����2PW�uD}�b9�����%PM���|�P~)x�?{���x.�Knq��u*K6H�q	k���AGҚJ<�(J�.ᬵy���,kM:�yzL͊�q���bF�����M���R��ӟ-��[7�d|���XP���|t�N�9���r�&U������G|M��[7�d|���XP����A�\�n���~�����G�٘�5߼
cަ��p�ϵ�DE1	�<������;�׊�:zL͊�q��UG�s���j�g��$Piq�VD�Lg�q��Dv;gJHn��z��r9�3���(�ʉ�I�,B�����B�[7�d|���XP���U8H�l����ײ]�4����=V8��H���o���&�t.�}w�n����|��T�.�l�.΍�7�"�����=���a�'�njVfV����x�%�$����{v��G�K$x/��&���7�ܥ��2�]Hf��?)�\�*�c�Uð�V���Z
�w�
8_�n�To�[r��}k:�(�U5ƚ��\�v��P���Ӫ��G�����x���`Π��yGb���u*K6HT�����N^!�"�{6N��p���
��|ſ��D�kt��9Wp��� ���U��7�ܥ��2�\Z�ؿH�jGjh�rO-�<i���A���U��7�ܥ��2�\Z�ؿH�jGjh�rO-�=|-�e1|E�A�2����ma��}.�����RE�s@�q��g�QX�QlxqG�T}�+a�C7�j��B���m l�o���ma��'f cTw��� +@����wF4��0[����	��N�Ae�#����ꀍ�����5	���]���>����C�h�'f RY%T��BPe.��xu	�>��l%i�-��9��稕�E����F��j��\w��0]ɍJ����j����tL��|g�Y�'���Xw�j�7��HaU$kX��a\Y���°��������ł�!r�dN�<@Iv��nt=:��(�
@��^y�~?�2vYl���#�]�!����M[��Ǣ+���G���"B��$I��w��,>����CΉ��S�|JY%T��BPe.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7T��a⨯/v�K7%'c��Et�p�VU��J)��� �e��uy��4��T�P�� ߌ���E����F7G#+�Ǘ0z�cUL�BJ��VR�^Ƒ����"X��[��Q[R�7��=m緒��J���W�7G#+�Ǘ0z�cUL�J=��'EّD ����R�^Ƒ����"X��[�'i�! ]���f�+��T���O'�lR�ܓ>��iכ���Mg)x�,��|��ZΫ��r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+�ڔ�wV���C�Sy6ג��̹��/R#�x���c=��V�j �F"������MJgrY��.!'Y��\�v�w�?�b�>޼�\�v�	�+�&I(&�L���mSP�]5����@�jO���a�pM�����!��"� +}Z�"��%o����?�}�	76�&�� Ӗ�tEA������L����Ҙ$7 �0��k{.Dt�0�Fc�9ٴqw_��>�ѻ�5����g�F.�u�?��'l���u�Ҷ�=SPn������`����8-|�D����<�.�%m�.�#7]��8���@�;����`Q0�j��9W����"�<��E�Vɹ���Ђ�Q�S���>�E�i�m}6O�D mWN\�.$�t �0��k{.Dt�0�Fc�{���"���@
H$��j�)�[���$���i�,�9��(�Ӳ�����±�sR�{F5Bn�LE=g��� ��"�8ߗ:w��Q/)�EY4d꽇��DlZ�G��յ[+8�^@Ȃ�z�wu����`�U�s��~-�S����"���v6"S���5i^����{ϧ��1���]��#�s���[�ُ��Ě���aT��3G6%�ȷ�F���`�j�{���"���@
H$��j
yd\V�4S�9躞0{v�c��Q��"��0����E�_������h�ӵeo�i� �x}��M����,��a9����vb�i0[����8|��]��0�ȍ�x�>c��O�"P���'8��)���"5�o٥yf�Kd+���A�,h�ѡ�@��6=3
���kd�$I��®�݅'�K�5ߧE4��T2����
,��y�c�M�`�TM�óM�˄NKYi�����.��B�M��:�گ��cB^�J*�Rs�0��7n������\�vŦݪ�h��-G���3��\�v�w�?�b�>��#�ڊ<?@���0���	_�>tt��n�{��l[hbvk~�#x��d2)#^`$�\����bs
a�=K�4t�4�;���Y��<�o��$��d�*��"~6���aq���`;m�!��nQ�rV���A�E������&<v�}��������@|������]�h�p���BHN��R���]�w%�o��]E����4|�N�f�0-=Y/�@��q�r����開 �R���d���M�Z�xuo��*Zx4���tŚA���ۖ�.Q�2�>�_����J�	�LÆ�[k�'��P�d�X�VM�����a�"}�=Ll���:���^�P�v�����"~6���aq��yx6�n)_�J�	�LÆ�:�;�������1;[lzRY�ȝQz(�)ةnQ�rV���A�E������&<v�}��������@|������]�h�p���BHN��R���]�w%�o񞾠����������3�RL�y�}Y-h��!��|K�{ߝA���:��% L����6���$J*�Rs�0��7n������\�vŦݪ�h��-G���3��\�v�w�?�b�>޼�\�v����0����KX��iknQ�rV���A�E�H/Q������-�z���3
�v�v-}�	mp=b�ɝ:�3GV���B�R���>_�?"������"KT���v�8:)��S��;���Nf�������M�W8�[L4���% L��Ȍ\����a���L����Ҙ$79=7��>W~4m�c},_⾊Bo�#���F�O��$�}$|~ïSup�xg쬉� }�=k�Rm���ӑ�xGe�;���N��}�!`���Nj�a=�S��j�����˓#���yB��K�Y۪	�}a�]�w%�o2�LpOJEl��Q�P�]zm?9ۄ&��%����"��y&I�3�b�}�IUr��Ӈih�|���he��G��֥��ع��F�9&t�A+gV���~�����.��4�F1��xs
�9tO�d�X�VM�����a�"�'n�^0o:���^�8�ʕ�Ke9Տ���i��q9�dԾ��?��B��]	�u�Q����������� ����H�ʱˡ�����Шr��_.�yE�ӜH�_0�g�ܧ�V*ڎ�0��D�9:��cSS�b�۪	�}a�]�w%�o&I�3�b�}�IUr��Ӈih�|���4 �DQ; Z�;�;}z&L!e1��bJ�5������қ�O��U���"�*�[�)�T���u�I�+�c��Uw���}�v���Lj��f=�2f�o��"��U�[в��*�p6�!"��֏����8!��vp�P}��O��^��mi9�g#����l���If�_���˱���v������*�%� �2S�;���;^H,�*}4��y������L�@��
<x\ċ�c�<U�X�HL�U��R8p��v;�}�i�pGա*�p6�!"tТ�1�y
���[�]��H(���Yy7uojr쇤���L}q��Ɖ���x ���r+�۪	�}a�����.ĳy�"�V��q&=�a�7�&�ҙ��C���}�v���Lj�󢘎��uҚ���"��yM�f�<�O���L��^I��'���: ��ao.\C�k���p4c����hl�6������1�R+-h]�D|�[�R"�R)�����J���6��� 8���;D��A���)x�?{��
0#`�1��JHn��z�6�����e�J�Pn\û�h�ם��M��_(����@҄���G�ۄe��D�#��%BJ�g
�zP�w:Ec�[�p(	��Q�^�y�zL͊�q��j.��?�Uʚ7�ܩc�r�(����.x�1�Yk�	�yOŮ���zAE>B��xf�� �+���/� �'n�^0o��N:�@?u ӫ/��m��8tȹH]g()��ikp���H���U�:�tw��΍�}����q�rX�]�)��0�E��zL͊�q���Z����p��R�}vJ^G�ɛ�!�~0��9EI����&��}����t����==�x�Y�E����F�_���˱���v�M}�nϺ����ڝ�ӡ���<K ���3�Һ�j_ R�ϱg#���
鴋��_�(�X�B;&��v0JHn��z���P��(��"�9-B���H��@!�#-�[ҭ�x��`��Ƈ_���˱���v��XҰ��
�we ��g�ɛ�m�d��b9���.M�"��Ӗ��ٟTP�u*ys!�`�(i3"�,�>E��ʆ�In��t{=J���y@����j5r�n0���� �}�jݭ�F����5��;y�O2뛨�2>�B�Q��>rM�Zc������3a���A�H�X����)ͶG�q�5իx`��:�T۳�͕���ȋX�b�t3B��*w�	�Z�X�ׁ��&J�b, ӫ/��m�h���Y�|ò���
��_�����v���-*���0i��¯�'Qd�i׏�����M\]YD�^�O�<om��Ts��E=����fU��b�TG|�wA���^�hŁw:����v�8:��J�m��iJIo�s��'��y[�@Ǻx�^�6/
�G!.��=x|]�m��|/���h��Jȶ�B��=}'t<��ġ��,�gXk���y�S}m� 2�k#ʘ4��\��sپ#�J��v�8:I�}-��^`�Ç(�/��@))�XDd�-$#�0$aX���ۖΜ(4���Yk˃TacX;���'?RgB�R���>_9g	���W���b���p��=�^����_T���a�aq�����x ��݉#���_J*�Rs�0�.{x>b���2��a!ֱk���p�G�ܢΜ(4��3�������acX;����*�t�J�1���{�H�a�\�#���F,�H��V�`n
V~$��$�J݃����t����~�/:��jsJ��U;���v�8:��jw����,�>2�0��&�)������Wz����vkN7pթ��ex�$���\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���И���ݥ�(��mK�cn��>8�2���H
.�oI����ġ��,B����s� J*�Rs�0}�g�*dǈ%�7:H� ӫ/��mO�%n�"�T۳�͕��w0H��G��9%2�8��!����&@��(+���<om��k%-uב8)x�?{��偗#���\h�x#�L_��$������Xjۙ�)��s���Џ�I��$��cn��>��[KxME��*�j�H��b�(� xܟ�,3JW̬���	p f�g�=�'��h��|=�^��զY�PG�(nQ�rV�)�YBa�g()��ikp���H���x��3�Y�^�х򪂱�j���Ү_s�=�����KC���x��N��\]YD�^�O�<om�����0M�C�T7���j5r�n0��:�_�B�T�;���N��6H*��l�A���ۖ!���6�,N|��|(F9%2�8����$}ům��KɑX�g���
�x��e�,d�z۪	�}a�iQ��ׇ��"~6���aq��yx6�n)_���fx'v�ao.\C�k�4yn���b�����V�I�e!��nH�W��3��oE�ƺ?Iߕ��1ҙt&H��V�K�1ҙt&H�#��3���׏�����Mă
�1��g()��ikp���H����-��԰�3�I))����A�m�(��:0>�ˇ̾\x#�d+'�tL���lϏt��B>�\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���LbFN��֬�lPCrM�Zc���o���Ȝ��(Q��;��b�=�*��i!�f��T1�"��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$��&��<+'�tL���lϏt��B>�\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���LbFN��֬�lPCrM�Zc���.�Q� ���(Q��;��b�=�z��Ce��f��T1�"��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$��&��<+'�tL���lϏ��E�_���\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���i�!�䒨H��@!�#-�[ҭ��F6q,/��h�`N���V�I�e!��nH�W�l,ѳ��=c�f������C;��?��QX��WG ����������we ��g�1P�n$~��7j�7'cT q��Ko.g()��ikp���H����-��԰�3�I))����A�m�(]�^Kҵo��(Q��;��b�=�v=]e�˽��q���3B��*w������ݡ��4z�Tqn�}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-���Y���� ��@s'R��E=���r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^��o�������|Iܲ��9m����uY�0��f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#L�tD:��@F�W�1'����
3����1�D�s &�`����w�ǻ��v�8:�^�U�3~�㕜��z ӫ/��m/���^��o�������|I��l�;?X�X��WG ���}��0:�{�.ᬵy���m/"�k�^��o�������|I{8��7�g()��ikp���H���X��WG ���D$��:��
3�t%9��s &�`����w�ǻ��v�8:�^�U�3~�㕜��z ӫ/��m/���^��o�������|I������X��WG ���}��0:�{�.ᬵy���m/"�k�^��o�������|I��p*_ �g()��ikp���H���MdGN����̾\x#�d+'�tL���lϏ���`3*�Z;�$ؔ�f���N|��|(F9%2�8�΁N#�ׄ��>��O˻����|I"n?��L�5��\�@���7�	j&f��w�'�̾\x#�d+'�tL���lϏ�B���l嬇uk���X9{lq�"�$��獶���_�(�X�f@i��������
�xL(�䆑�֬�lPCrM�Zc��_�-��1��r�.Gb�TG|�w�bX�T���5��\�@���7�	j&f��w�'�we��3��we ��g�1P�n$~����A<=ж��˓#��͢��V0\�Q�%,��7n��I+ɦ۫K���L���4�04�jfx(�i��/R��!�ˢ4�04�jf#��`*;T�g#�ˎ]":V��ak�m/��m����e�,Ÿ��U���:k�ף���l�����;�R�I͗�ၚI���ln�λ�����E˷\�H��/SggR��N�$���\�v���K�P�%�Uʚ7�ܩc�r�(���JHn��z�r��]�]��eCǮ��\�v�JE|Q�R�hbvk~�#x���EE��&�FO�r�&U������G|M��b9���M��A���va�{����2����%��/q|Ld�r:ha3B��*w�B4~��	��b9���2s��f��6������1�R+-h]��857���Ѹ�*��7�?	�^�F���.ᬵy��ҀD�C�3'�a�e�7�!-`���wԸI))����A�m�(� 9':�&'��v�8:��MWU�?
�%��/q|b�����V�I�e!��nH�W��b9����2�u|���U��+�X��ѐ$�؞�v�h�Ů���zB�$�yRGy�ˆn����N��+�[�{�M�>�'n�^0o�!O*�]�۝,E�?����S����)x�?{��{P���J�	�LÆ�(�.���{=J�������e�gb�TG|�wA���^�Q�^�y�N��B�)Y�+U�HJ�hY���ZSu(�Y�^��	'gx�u�%Ah�%4
>�(_�<�� ��&IWN(����l�����r�3�����!%Ah�%4
>��XP��ș�_T���a�aq�����x ��݉#���_J*�Rs�0�.{x>b���2��a!ֱk���p�G�ܢΜ(4��3�������acX;����*�t��+U�HJ�h���)Q���3D�� <� �|��� �b9�����6*�U��'��pmp���s�&
��3D�� <�7ć���l0��F��jȨ�� "���!h�b�TG|�w!���+���� 2�k#vO�1YK�8���l����׈�	�Ȟ�����hLKW"�,�>E����\�vż�ߞ�Kе�B7S��A���9!���M�V��[� ӫ/��m}�g�ޢ!6������1�R+-h]d���85��"5�o٥RK܃��hbvk~�#xz�Ŕl������k!�tt��qN�����v�0��YB��F܂d�ۤ�|��F�� ���3�Һ�j_ R�ϱg#���C�'���#�A�6x��+���/� �_���˱���v�0���f70���!�`�(i3 ���3�Һ�j_ R�ϱg#���I}��NV�MO���9�<�!8	�I]��� N��r*�$��ûX��kRCլ�����`��&f��w�'�?t�kJ �&{�zYa���<��ɢ�U8��ّ�k���H��@!�#-�[ҭ�g���y��b��v݋N��������c��>z�Vg.N�������6���|��"5�o٥۪	�}a�iQ��ׇJ�	�LÆ��/�i�����܍w�S}9g	���W���b���p��=�^���3
�v�v-}�	mp�����2x�N?Dd�-$#�0$�.�-v�Μ(4���Yk˃Tc�δ�0���'?Rg�\�G���nQ�rV���1���X��WG ��D����jF��b�(� �	T�����3
�v�v-}�	mp�cA�N�Y�74��LM�(�� 	l��lBýO����ezꥦ��r���:�����C��괽���5%�"|R��9%2�8���x�Y�1G�Sזi�)x�?{����ҳ�ET��o*|�[3�^�P�qjhbvk~�#xe�����t���3��Μ(4��fU��S��ɻ�7��M����v�l5��� rư1�l�_�4��׏�����M\]YD�^�O�<om��Ts��E=�!�Wƞ$�FA��mӡ���<K�hŁw:����v�8:��jw��.i:�����n�{��l[hbvk~�#x��d2)#^&|���BY��l��=5;� Bw��A]k �}�Y�PX�)��s����,�Ğ<�q�;���N�?~h��dg()��ikp���H�������K%��C�<GUl��P��3�(��mK�cn��>8�2���H�?WY��c�#���F{\��@�����p��}��aq���3�ãK� ׏�����M�8�� ɮ�_�(�X�<�q��Dp���$�J݃����t���Ԓ;7rgb�TG|�wA���^����}��th�U�CLf�� ��nE�g%�?Iߕ��1ҙt&H!F�Mub��ġ��,'5��'Xhbvk~�#x�o���#�51��r�.Gb�TG|�wc�'6���7�b^��!{lt�m�����ݟ���O�͛PA,q �?�2R��b�����V�I�e!��nH�W�yl~"�u]�%,��7n�W�{�'�h�����	�����A�\>W�/Z��B���[@���[��QPw��r|��߇(������x#��y1jU�$[���
�x��z�?<t��s��U;4�a&�bB�i2n_����~�/:��Ż�&ǥ��a���F4�04�jf���w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m/��������|O�\�+�q�� 6x�@Ts��E=��T7���j5r�n0��23��-��2j5r�n0���Z7£�&�x(�i��/R̬���	p}��%%��(K;�I�N���	>����E��Z���HB8�	S�1|��[��H~n�+�W�z|:)��;z1
8��h.�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��Sa�4o�̽��h�`N���V�I�e!��nH�W�l,ѳ��=c�f������C;��?��QX��WG �����w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x������|O�\�+�q�� 6x�@�����3��#�[��T�s Wd2uUrG���L�͛L�_�n�To�[��g���a��>�8-�ށ���
3�-�f.�o>��O˻����|I����ZqM<O16�,��p���#4�Te͉�Xk<�zPӹ�&���Q����N�������_�$��o���*ٝ�/�K^b�;��	+�uG���=���[f�[q�g���!_Ez�1[FQ������-Kff���e�F�N�@E�V)�jP|B�1��URpL���q���3B��*w��&�Fc?�}c���x��z��d>Q���G&o6_��'����Kf
�f�3
�v�v-}�	mpҭ���^���b��v݋N��������;B�駮h�`N���V�I�e!��nH�W�l,ѳ��=c�f������C;��?��QX��WG ��\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[��m��I���f������C;6�GRe��X��WG ��"�!�RMUt��!
*J�K�b��v݋N������&I�~Wm@ˎ]":VȠ຀�m@,5��*#y֬�lPCrM�Zc��s�I�A螗|�S�
���N�@E�V)�jP|B�1����}�\�T�s Wd2uUrG��÷=%s��Gy�ˆn����N��+����x]Q*P�#�f�D��&{�zYa�9�LL;M���7=�[G��"xC��-�T(u	M^��|A�Iu*�����4^i�u�J*�Rs�0]�����sk�����\�H��/Sgf����O�9<~�p_�X����)ͶG�q�5��5v؊	�\�G���nQ�rV׃_
"Y9<~�p_�X����)ͶG�q�5�D������aq���5�*��֕�T��̪mMUt��!b�4=y�(ͻ� ���7���ìL��-)6������_�(�X�f@i��������
�x�<zf�L��H��@!�#-�[ҭ���;v�H.h�o���*ٝ�/�K^b�;��	+���$!�+]�4"��B�*�A���ۖ��Rg�3e�C*y=�_�n�To�[w��{Q����$,��F܂d�ۤ�s�����z�F���D��݌ߛ�#���F,�H��V�`���$,��F܂d�ۤ�s������3
�v�v-}�	mp<A��^\[�Q�=ؗ���`;�nQ��A@��sZ��o���*ٝ�/�K^b�;��	+ѺA�⿷�3D�� <@��fG�3
�v�v-}�	mp� J�H�ޭ�2�q�]�>��O˻����|I�w�63xHl��7=�[G��"xC��-�T(u	M^��|A�I֣8kI�g�I))����A�m�(i��C֤�we ��g�R̫���+w`�M�F��H��@!�#-�[ҭ��<���\Q�b��v݋N������L�{���\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���Г�D�i�^�Ax�`Vk���|�i�!�䒨H��@!�#-�[ҭ������̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-��|��������2���t����)L��b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tF�W�1'����
3�м�1#���q���3B��*w�eB�_f�f��T1�"��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$c��X	��MUt��!v6�RMS���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��N���8@�we ��g�n�J+s����$,��F܂d�ۤ�m�>!������ᇱ�����s�`�|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*;̊���z�1[FQ������-K+�0�xT�5T q��Ko.g()��ikp���H����-��԰�3�I))����A�m�(�A��PmP	�Ȟ�����hLKWਠ9V�-^֬�lPCrM�Zc�󲄊�](x�%�(^?�f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#L�tD:��@�JﾥI��P3�lWD˅yw���-u������b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tF�W�1'����
3=�ЩT�63�q���3B��*w�eB�_f��0?2�U�w��r|��߇(���л���.Ȃb�����V�I�e!��nH�W�t<wN����#��%�T�s Wd2uUrG��U{��b$v��`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B���Y���� ��@s'R�.R��д=|��(Q��;��b�=暚cpSi�}�vo;��|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*;̊���z�1[FQ������-K��+�v�zT q��Ko.g()��ikp���H����-��԰�3�I))����A�m�(�A��PmP	�Ȟ�����hLKWQ�@&�?�֬�lPCrM�Zc�󲄊�](xDe��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�X������<�N�����K������:^��2I=����P�7n�+�9�#�PA��n�{��l[hbvk~�#x��d2)#^&|���BY��l��=5;�D�A�'�Go��<e�Y��%,��7n��A�N�'�]s������&{�zYa�8��V�嬱�4z�Tqn�}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-��|��������2���t�h�N#�Ǐ��˓#���6��R��O+'�tL���TĆ�AUt�\�|��������2���tԷ���t���3D�� <�1��h>߉�(Q��;��b�=�U3{����B�L�͛L�_�n�To�[��Oy�,��a�z6�F�W�1'����
3Ts��E=�L���1;Lxz�1[FQ������-KǷUv��9%2�8���A�+���i2n_���Ŵ��`���H��@!�#-�[ҭ�*=�u�8����ڝ��Ҟ�T��7}�t�ё�F�]	
~ao.\C�k�Eg����0˞����Ti�^�Ax�`Vk���|�"�ϴBꙕ�T��̪mMUt��!.���9fj�}�Y�PX�)��s���}H]�˖��1ҙt&H��I����8�����|I]��ם�y��1����Y�^���Y��H"��h�e��SV�$#��Dq;��*�\G�I))����A�m�(�NjX�U�4�04�jf�5ߧE4��k.�C��(~�;���R�`;�nQ�Ǡ%"t��\�.$�t�:����RW@�S��o�C�ޝ9IR���c&;�L�FZ�1Ǩ�Yc�A�/����<.+6J!�5����`Kְ�4'N5wĒ����H���o��qo�:���$��Xo���~��1�51	�<�����ȳ�%�MZẶ��Ϊ������1�/؞�{�����eD������~�7P��T���\�vś��Z1`� k�|6�8�\1�p���j�L��G�Ӿ�@��[p8�]�1d$o�[\"+<�}��|~9:6D�� ��;J�o��]�����G���K�*�7`����M�Z���	���}0x�5�Y�w���8���N�:�eEJV�����a��&���O��*�����2+C�	�p;�j�`,k����}���Br���l�*y=�8�4�dL��p'Ik��M�Đm�L��X��O�J�t���V�����aǯ�sE���yL6C\TF��I��RhF��C뻁�ih`�ol�Ǯ�����4�k��Ȳ2�Ԟ-zq��D�	a�]a��1qh_�n�To�[�C��-��JHn��z�Lqܳ<��J*�Rs�08�b(��+�w]�B׿�ġ��,��ȧ�!^�x���\�2
��F�l��=5;GZEh5���'n�^0o��N:�@?u ӫ/��m��?�4D+V���"�V]a��1qh�>z�Vg.N�����[���S��IÙ=�H�+������eiVc�$J�{�����~�Bhl5�v��fx'v�ao.\C�k�ru1�(<�!ֱk���pF��kL��r����%;�%��/q|Ld�r:ha3B��*w�B4~��	��b9���2s��f��6������1�R+-h]�+� �J�����0i����N|��4���ߗ6s�B��@N�柇���j����rN�ǁ�f�T=�����JHn��z�F�x�aK�k����k!�\Z��K��ϱU$��0��иܖ��R�7��4�����I0���ԏ�.fOe	
���}L)��b�7�/���^�cm��3\ql0��F��j�
����uK�I4��欱���j����S��3mU�r��>'���}�pIɽ�Jz_�"�,�>E����\�v��u����)����k!�\Z��K����"4_��%��/q|ܴ8`���r%��ɷ�C8��+Z%Ah�%4
>��XP���a��+�R��$:N��ܙw�F��)�j�F2I��'�(��_�8)$���}6=(��B���~���}�=Ll���<2
��ױ��.��B�M��:�گ��cB^�J*�Rs�08�b(���os0c��ZLN�	��`h�-�����0_hW�D$2���O9Կ�eJ}v��.�x z�Jm]A�/��� �R���d���M�Z�xuo��*Zx4���tŚA���ۖ�bݭ��s�J�	�LÆ��E� )�&V���"�V�p-�8m���DŤ���uXSr���K�H~S{xv�NI�����G�	�Q�4�L �׭t��y(���F�
�UE/u����`�1�aw���q���0/�Ů���z�f
�u��4���Fr�g��� ��"�F�*���_x�]�V����ߞ�K�o4 l�5Y�0`�WC����B{�LϬj�iM�!��i��Nc>�V��v�'���Q��K�Z�b8�1-�ĩkG�Hl�W�uXSr���K�H~S{xv����K8 t����%#�����m�%f�QaK��hW�D$2���O9Կ��w��E��0Ů���z�6o[��:�-$�I����Q��Ka�gN�3cx�]�V����ߞ�K�o4 l�5Y�0`�WC����B{�LϬ9{vw��~�=D���C�9Wp��� ���U���Q���(�r��VYW\�o���*ٝ�/�K^b�;��	+����4���XP���3Zk�E��% ��q ���h�c�M���v�8:U��z��!�nQ�rV",�Ű�/؞�{��X�i�R�ռƐo�c�?EcD�=1]�Ed|�+���\�vż�ߞ�K�9=7��>W~4m�c},_⾊Bo�#���F��-��j����猵D��I��'�����7���{r�����ތ�1��\�v��\aьIR=Ϊ�/-T)x�?{���x.�Knq	6�q�i�d�<om����t��W2�A�;�֋`NY~�y����u{ᵿ����KƠQ/Ǔ�;�CSW JI��'�����7���{r��f���꜅�R��ӟ-�1#��Z�����XP�����w�K�b��2W hbvk~�#xǩ"�4s2nQ�rV",�Ű�7���8����v�+ʢG&q^�`
�c��><�$�X~��\��|�^��
�>IÙ=�Hss2����`�|��K�z�H�MPq6.?�)���؀qjZ�`�|��K�z��|����=%+]Bo�A;h�F��O�i���AԢ�a\�D�����R�`�|��K�z���k��$a(􆿳����d7\�{"j��?�o>����h�9��c_����+#��.X���*"v%)��Qcm hP"G�wk��r)��ׁ�a\Y����)���8˩��F�{a(􆿳��?ƾ�؀qjZ���A3�(N��㎏qló��|�����V��ߝD9�{��灊�O�i���Z鎬�������(���`$�P.eE���lC��U�T�\ ��y�.�`L�P7koеI͢'�����t$I+�V�6IWJE�YY���F;�I�e�,��[�9q�Y�{'%s�h�v��T�v��1���6��	���`y���/��=6�s���l�%��iA����
_�n�@/%{�;���$H<�7̈�A3�(N��㎏qló�Q���l�G�p�PH�^=�h{&����������$�1��i���E�ۡs���ψ�A3�(N��㎏qló��|����=%+]Bo�A;h�F�`�"Q��:�kw�j��-}�"��{<I@1��+d68&~��0w�y]����^��t�������QOm��/a��\�vŶ�T���R�^Ƒ����9�m�~��#I�90gA�I�y�?ܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'��!�a�~s����R9Y�}��`y��� D�f'�o!�gsM纞��G�٘�{����#�r�s��l�dט�w���f�ܗ��DX<�c>1K �:;k�+��b9������|L�K�)x�?{���x.�Knq	6�q�i�d�<om��'@�(��P�����k!� �J��/�oxW�}�zX<�c>1K �:;k�+��P4ǲ ��V �-�{q�������ތ�1��\�v�M��r�&�(vW4��`��?B��ž�'�t_� �e����Eck[�x�X��u�?�=�r�@^7&ģM�'n�^0o�<:�W�_�l�J;�RQ�y�� Y{q����'6���;8=�g��U-�e���TL�b�������z��d>����C����ud�Ad�'n�^0o**�ХM
��\���ǖ��;^�6#9���k��$����y
��J���e͉�Xk=��t�(�e�;����J>п�p=	�˳͠m�xW��9u$d9�ל �w.���/�K^b�$����oh`��E�hxǉ �Ş(�/�K^b����RXĨ�z=R\�U_�+X��-�&a)��V�t`u�`�|��K�z���k��$����y
��J���e͉�Xk�
̄?�9;��0����GI$��ǂcY�~�s<��MRZ�α]�H��7���ìC������*�H`�~��ƴ���(�_�8���< �w�?��ǉ �Ş(�/�K^b��6&��^�<%̚K"��+Bo�A;h�F�����`̢bޡ�W/S��8(�E���Kt�5c������\7vm�܉��J���e͉�Xk/[�^��`^r�m�����ч��,1��;p���#4�Te͉�XkN��"�&CA��E�9<Q|Z�j��?�N�@E�V��Ù���_�n�To�[_��ƕW��Ĩ�z=R\�U_�+X��"M�<	I0���ԏ�.fOe	2S�İ��y�ѱ.��tGy�ˆn����2�-���J*�Rs�0:`D�h�#�*"v%)��2������3
�v�v-}�	mp��8#�&��Y=�ĵ�"xC����=N���#���F���.;����\�v�g�W�I�@T��*T��<om���}�և^H��/1A출�k��T9s*��ԜF�����t
��P"G�wk�١��	;q�J�� m�h�5,Wlr�r%)cA�z���a�R�wX�Ց�~�������`~�ߪ ��e��R��!kr��N�؆�B��W+`�x�oP��@t�&�e�5
��x4ca&	���Δ���7�j2�ٯ�e������sC�|����1�Z���=�Ln��S�W�כJϾ�i�I7��-5r����%c��P=@��������$��Xo�U)+N��C
2��Ln��S�W�
����uK�r�&U������G|M�y+�>K�V,�v����f������C;��S���'n�^0o4��t-s�C
2��&~�� 
iEE�Gp\匔'���� ����H�ʱˡgb'e�W�'n�^0o�!F�;^/K��^̽1���C�M$�;5M��)�$�+�,MN���OON�
_�n�@/%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7���i�_:�����k��$a(􆿳���L��F[Ԃj(��VX����nU,�a�r����Eyp	�!�*��2}���5�Y�w��qsd���Z
�B�uJL�k�Լ&��PW3��P��/؞�{�����Go2W��,8����;A3�@�����tS����'n�^0oˇ��_S���$:N��@�1�˓�����f�l��=5;$]��Af��v�c��Q��"��0�
MQ9�F�����
��\�H��/Sg�w��'o�V���"�V���Q�9e�۪o�y)	�'��ɡ��F}�$xd<��\�vŊoC����$\�H��/Sg�w��'o��ڎ5�����>z�Vg.N�����B�L�[��OY����A�b��v݋N�������`Q�>=����V�X����A.�%A��C1#��Z�����XP���	3i�\��׹��t˻�� �
n���@q����Ǎ��mjR}�����S���'n�^0o4��t-s�e0��Tqmp�AJ�e�$���U�D3�f�Nd+l�t���c����f�����eR�ʨ��_�\G�k�y'��aLn��S�W#w���	(���B���Q��ǺΕ�V�܄WD��|������F�QY���=�w�Ηե>���Q=z����9�r�)۬
Yz,�o�oF�����ư�h-�j�� r�[WQ�z�וy�+"�)lCN��Ҧi)D��%��Q�R�G�)q�j��U�T�v���*T�@�sJ�|���"��|���it	�TU����z~[x�h�E������x�@eӎ��^S�^%��&�I��������"H��l%BjW��5�A� �cۀ��%a<��A.l��0s1i�f����0+W���F�^�Y�7#�xI���|�r�HzL͊�q��/�"�=bߣ$5/H�<u���(�?���it	�T$x�����7���8��� B^�.�ߘ�)�I0M�/�s���'n�^0oPpkiq�o�H�MPq6.���fa���ӵ#yӛp�Tr�j.`#2��%0d�.$s����c�w�i���+�r�2�=l(	/K�^0N�mC}���������I���9�"E&��� �Z��T��B'$��k��P=jǳh�5,Wlr�r%)cA���ˎV�I��'�Q�%�+2�0M�/�s���'n�^0oL��w���GF��a�1�Z���=�g�R�:M�BvGޣkQ�A���ۖ�k�V\��P4ǲ �����zPuZ�v|��3�%x��GD@�F��q��W�����לo�	�r8S���Qi�4umJ:%�b9�����%PM�V���"�V%$qr��pa�Y%�^1#��Z�����XP���G�@[E�Bn�*5H8P�x/���������ׄ�Q�K��t(��u��n�{���G�ܞo�$C�p�AJ�e�$) u3��`��U��.м�\�v�n��l���&��K���E4J�VB���;��%YՏ���i��*����{�"��}�
�'�!�K�|q��=H��6�����рӚx�2�V�aֺ����zP"�k��ir'�yK�w��b9������sh�f�)��u3|ڛuC,h�Ʊ�_�eD�I�:O0�9C��d
���u[#�g�+��8�΋�)�Օ��qvdЧ^{�jX�#���s�6�U�D?����M�;�>���1p��N�oJ��JHn��z��S3W�K@S������H�|�ߦ��X�G[�Q��ǺΕ������5�3
�v�v-}�	mpŴY����;���NA��sm.�9I��'�N6����(�;UW�������4���XP��ȫ,Ÿ��U���:k4�9��S�b��v݋N������oV��'wNF:����Į��KH ��*PX�KL7��Ѹ��R["��J*�Rs�08�b(���zY�l��R�}vJ^�?�1�{Ů���z[R�{ EE����u��h,%I��t�'n�^0o<2
�����L;ø\����?v��0\�^�� ӫ/��m�,�XM��v�c��Q��"��0�z�qw ʲ��h�ӵeo?��`�1M�3
�v�v-}�	mp�i��,zx�����k!�\Z��K���8մ�6B�ʻ��AN�It�Ɍ+8�3��$<�Q�R�j�`��2�.�05k
��F�2�q#O��*V<�ɔ�,���T�K�TZLk]�V�Y�\Jm�A���(���d0J�̛�ĭms)������*��?���-)zd70ǰ�5aj�r�[�"�@��e���ú��'��X�T��A���sG�]b�` ���"�+�*�p�a=}���dm���lD��~��~�
�t7������U�M��	[�/��8!�`�(i3зq8�Ј'���Xw�%G��ly�Ed��>�^���n���g!�`�(i3зq8�Ј'���Xw�j�7����`�z��Y��)�k�������x|qj0�vے�(�iF��׿]�/�˟��7<���������	N^�U{xN��i>r�<Uee��~j�j����.��@����gGKCYb,�q@9
!�gwe�ŉm�m�jp=�>��o�
�v�ξ���Ix���Ka4ؿ�v�ct�:��RE�QS����>��"X��[��Q[R�75�e`��9��əS\�
���X��d�٣���������ݹ�0���f�Nd+l�Yҽ֗�?��}�ͭ��I7��-5��6��	���`y����@����gGKCYb,�q�U�`��dgwe�ŉm�m�jp=�>��o�
�v�ξ���I��RhF��!{X��U�B�ʙ@E>*;�¬pX��g��U-�e5��e6²�23
����X%�(���z�w�s0�W9a!@�'b�t	�U���C��O]r�<Uee�N�����z%$��h
P�%.^F�	��lC��U�T�\ ��Z��| �Ɛ����n9�}��������-�`~ ����i�0�OgA�I�y�?ܔp�l
d�R�.��On��M���o�G�m�?H�OM��`�@����gG_$Mt�z�N�X�!K9�:�a��Y�{'%s�[�&B�踫g(�r�x�y�Zgl,�B۸��ʙ@E>*���ls�u°������R�wX�ո@����gG�T8�����_��<덲��+�J��Y�{'%s�[�&B�踫g(�r�x�y�Zgl,�B۸��NI�:7�N�5�%]���a(􆿳���2����.)}���/�;���_!�`�(i3	r�&B"K�͢'����&���Z02��`�z����k!�\Z��K��ԒZ	x�B� Ei�lmZxE���8��?��Q����]�!��	Ǹ�y85�����5��d5�:�w�+���LQ���"X��[�z�C���|�F7�_����dn��Azg���d�٣��c�A�L'��Gr_���GF��a�1�Z���=��L;Л�����Øf}�
�?��h��=;���,�Q�'���Xw�j�7��Q�%�+2�ƃ
ᾆ�x�T�\ ��i3�|)sՀ@�g}��c��lmR�S{}�d�٣���N N�S�WT� �`�o�:���f���Iv)`ɋ�ġC���}�
�?��YN
��)ee���b��U,�(�)8���0y�	 ���t��h�/a�'�̗�����C�M�����T�\ ���|.�Tӏ�;��[TM��a�D��<~lf�;��z�f���,(���B���̴_��EI?�R��n��am�Za(􆿳���Qs���Ѕ�HN9�âq�t�d� ��^�:AԢ�a\��F�dH�Dj���G�Օ��qvdЧ^{�j����#oM|#9���b!��u��4br��BڴQ��q��T�ٮ|�,
������|�FIsŭf�ҿG�p�PR��{�&�8���/�a'�<� \f���ѩj��Q?r]�������"����Δ���7�j2������%G�{lGD�V�B���q5�n-�@�4ڧ��~��r�pzl��a��YN
��)es��S������x�@��*��1�G�p�P�㎏qló2u?r���Y�G�˱�ߓC娤l����0"yI1/h�5�G�G�d�@���Gғ�vq�\[$Q��
�̞��>�nQ�rV�}!�@�?0a(􆿳���Qs����p+�@���5���u�L��E����F��"xC����=N���#���F޷�����j�׎o�|��he��F��"k��d�o/�d��7���ìk���͖w7a&r"� L,|��{>��Rr�@r/u���� Ev���J���e͉�Xk�3
�v�v㍼�@��⇋g�DE'���c�e�B��G��ӗ2}�<��b��OFJ> ӫ/��m�y:�u�Jq���wSK�T:���V��pu7����d�٣��c�A�L'��!�a��5�%]���a(􆿳���2����.��DP֞ cVe�U2�<�n`5�fK��0z�cUL�8� �,������]'m���G�K$xE�p4rqG7)T&I2WM�R�wX��}�
�?��ƿ�d���зq8�Ј'���Xw�Y�r�7"�[�=�5x��A~*aiqq��T���E@~����`y����@����gG��5�!�m��E����FZ鎬������_�,�;�7���c��չ�Ad��d�٣���N N�S�qg2�K?\K���~N|�H>+�w�\w��0]b!��u�#� �,Wɒ��r����q���U��@����gG�?#dK1"�`�	���������S8��$FW �9�װ?�p���5�%]���a(􆿳�$��ı�o�7��"=��G�3�p�\��C,�2�!�`�(i3ғ�vq��/��j�3�T�\ ���ό�]2〧I���/s�1��p��lJ��튝�b�Bϱ���w�K�b��2W hbvk~�#xTU]O�d��g��U-�e�n�r{g�〧I���}�Z'BY��lJ��튝�b�Bϱ�a(􆿳����^�򯊁�i���,v���p�m~|���A�X�w�?ׄ/�L�^�Q[M��&d�X0��±�sR�{F;�f��X���n���k���#��(����@Pe�?�@��O���d.���}j�>�`htu�Ŗ6$\Kʍ2ӆ	+��[X-�BM�ܤm|��Z�j-J���\�vź�^Dv�7����0/ܤ�(g��V아�nu�����.>mǐ�? J*�Rs�08�b(��n�� ���'�̗����#!d�+I0���ԏ�.fOe	��Cja����.)۞O��\�H��/Sg�w��'o�;��ވ�H��=#+��^n�r���n�(D�G�\ϫ\ʃ�1�9M��p����=j����s̓O "*B�^�b\��{��7���	(k�t �j�&.U}��le5�`���pɷ)A���	��s~d+�T�֓S$Y��C�9I��@��F��6�y��Fp����f���,(���B��\���V#��p~z�r,�b��r�
R�wX���7�b����'���+)'J���|�b1�#��d_xZ��j�
�iB{�Z�_��?� Zh�R?�R��nI4�p� ^�b��v݋N�����~DJ��/�a(􆿳����d/h�5�G�G��*�Աߛ+����m�W�h��8�
,FI��{�F�S��\��g�_2���� ���c��(r�x�mC�n[�=�5x��j|�>�Oy7�x�����*ܑe�W����n�4�`t��D����M����A�m�(��ڽQ���}�
�?����'�u��TʯF��zk�:A�	S�r��AR1<��J�@Ym��`�z��Y��)�k������Pv��On�T:���V�����,Ǣ
��p��媀?��(��I@1���t$I+��f�kN�ı*�7`����M�Z���	ԒZ	x�B[�=�5x��M��%LS��b���jp�B�E`^n�&�
_�n�@/%{�;���$��dg0J�I4��欱���j����`t��S��K�Q�3R�e��Ӵ�"�6j��;٬sf.�@O;^p�]�|��{�r�]#I�P�*�7`����M�Z���	��"X��[�z�C������N���c�v�J��sr�l�k]m��FAN���d?�o>�R��}���N�ǁ�f�T��p_U
#�g��U-�e5��e6²]�N��&���3�L���'s{	�h�v1a{J�;J�F�`�|��K�z�Q���l�N�����:��6}���8���/�a'�<� \�U&�Pֻ�I���I���C1zh�,0 ������c�SD釛-���>Tf�Nd+l�Yҽ֗�°������R�wX����K�Q6��~p�=�J����6x�F�-t�\��ot��c�SD釛-���>T�=�	o #���}�pIɽ�Jz_��|.�Tӏ�M�]x���'b�'=�(�ժ�E�$��*�]u�l|M��?T�a\Y���{lGD�V�B	3i�\��׹��t�'jG+�$�H���N�[�s���_����J����]f�*Ƶ �d�٣��c�A�L'�d;�T�1�a-���7a
��r�k�Ղ����Y-��V��k�	�"����G5������
�CӞD
ɴ��z�D-'��7�q�����,ꩊ�q��T��J�s���
�k��!a�tc�&ck��Wڭ��h�Ɛo�c�?EcD�=1]������R�wX����K�Qɲ�cz���ł)w���m�±��m|�0�n�6J1��J���e͉�Xk�]?w�U�]��K�Qɲ�cz���Ӵ�"�6j��;٬sf.�����ֿ�d�٣��c�A�L'�d;�T�1�a-���7a
��r�k�Ղ����Y-��V��k�	�"����G5������
�CӞD
ɴ��z�4�	���WdM4@��B?����P"G�wk��r)��ׁ�a\Y����+���LQ���ll��4�(�hF�w���a\Y���(Q6D����z�C������N�[�s���J��sr�l�k]m��WD �6�\5Gy�ˆn����N��+�29
����
�CӞD��gn�=4�4�	���WdM4@�{0	�b<h� X���/�K^b�����4��g/�Q`���$���^��y6�T���1���;�{1��]�N��&���3�L���'s{	�h�v1a{J���ӹa��	��"xC��}Vq$GѲ��W��mTS{lGD�V�B	3i�\��׹��t�'jG+�$�H���N���c�v�J��sr�l�k]m����B�B碕d�o/�d��7���ì�"����x,����aR��n�J>|�
#�`�^{��u�oD�|.�Tӏ~�L���vi��N�N-��;��M�z$��PЧ0���ö�z��d>3EKrM3�Vy�oY�E@2u?r���Y�G�˱�ߓC娤l��3>�3ʸNݓ��E�/�������� �mDƇBHx\�'���Xw s4S�'�i��`�z����k!�\Z��K��(Ko�yؿ;-;*�7��;mQ��8���/����,DTc�~y��i�v1a{J��H����� �����p՚��l��Hr�<Uee���R�}vJ^�k��76���>k��@����Y�Ө�՜w��yy����i���~�F#3���T�٥��T����P�H�.|�eHg�w?�#�h&
Qno��9�?�6��3k�勿���L���N�b�'Be�X�;�Q��[<!��e��N�@E�V!:忴�n$��O�&��2�0�5��Ɛg)x�D�����X�;�{1�牽Oi9L�:�k]m��|m�	Ƙ�z��d>����C���cׇX՟���K�QR�Xe����ɲ�cz����n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7����������n9�����[m�ɲ�cz���7s�9���o��S8�/ #O�)R�^Ƒ����"X��[�z�C�����DP֞ U�����L�����eK媀?��(��I@1�ؠ&���Z02�=�	o #���}�pIɽ�Jz_��|.�TӏU�m#j[��i��z�d�����YDl�L��M�,���	N^�U{xN��i>�/�n>�.-,��Sq'��_�H����K�Q�L�t��n#�%��>�;����K~���A3�(N��㎏qló2u?r���Y�G�˱�ߓC娤l���Mq&����	�A��ԡ�f�s�G��3�X&���g�<�>�ݙ�1|�דu���y=� �e��
_�n�@/%{�;���2�0�5��Ɛg)x�D�����X��9���t�����_zx��@S�@��NX�c`o�Z鎬�������(����}�O����z�C��Э��_zx��@S�@��NX��gﭔZ鎬�������(����}�O����z�C��ЁZ��[s�ǖ��`Y��E����FZ鎬�������(���SG㴊�?����q5�n�JrPQV�R�wX����K�Q��6U(�<",�Xʚ@h�d�٣��c�A�L'u�6949%t��R̕q���s���8���/�O�&�����)������F�O�_եS��Q]� _ό���.���K�Q��C�_���O؏����:7s�9���oC�M��N�ہZ��[s�{���`7s�9���o��S8��/�Vv���$:N�uWX@z�(�%�8���Qs���Ф��=�W�ۻ�F'i0�UF�o�$�d�٣��c�A�L'u�6949%t��R̕q���s���8���/�a'�<� \�����5_�(=�oaJ7s�9���oC�M��N�ۭ��_zx��*%΢Ӟe�H5��M�0�W9a!@Q2�+�Yɠ�B�D�F ��hi�aDU�G�a�E���Q]� _�rs�i��d�	�6%m���������qW[����Q��Y����Qs������b~��L_��f��<<��%�7s�9���o��S8��A��H�cB�pa�Y%�^(Q6D����z�C����S{�-CK)�yy ={�%���n`5�fK��0z�cUL��_��h��Jc'�yK�w��g��U-�e5��e6²�[��s�a0��#�����\t�c+��d�٣�����6>���ÕB\�6NtNF5��q䆆�$�\��i�#�:Q2�+�Y�'@(s��k����PĐ�ð?����UЮql�N� �$�6ֆ �Y�ƽ���j׳�)N�^1��.�B�n&?�qi�����f�,��o�k����P��)YL9~�Y�ƽ���j׳�)N�^1��$��劆g���!a�`:O�����I���Z�΅��u�H�IP�,�o�*$�n��,�Y�����|�å���inw�T�yp��&M���RV�h�6a���y�X�,4�?nO�J�t���&��}�b=�Ea�\�+���wy��urY�Y�:A0�,�`�_������6vV3��.@�k��m%	' ��a�I�..��/��ˉ�c�}�C�-�X]t$I��2�b=�D���u�\ssf<6A�t	�a�4)�k��D9�$n�0 *Pv!��\�� ��z*K��I4��欱���j����|�厡��� ���y�O�W,�P �P���UX�� ���JH����8��#I�ND�s���H�V��^�5G�����&�@�}�-��w��k]m��p�Ńۗ}:�,\���ӟ�X���&�@�}�-��w��k]m��;����)�#qp���W/S��8(�E���Kt�n ~���7��3R�e��Ӵ�"�6j��;٬sf.�5^����r�^E4+у��b�Bϱ��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$����Od-@��F~*7���&�_$� %7䨁c����t& ��i�߬�F�<|Mabi�~�-���G$��P���UX�� ���JH����8����F)�~����H�V��^�5G�����&�@�}�-��w��k]m��p�Ńۗ}:�YN
��)es��S���.�<Mm1���P�|T����E�E��3�L���'s{	�h�v1a{J�d�	@f�u �U�N;k��!a�tc�&ck��Nx�P��A���TaZ/����>��i��N�Na����g=E�g�N��S�yN4�S���%��N[�[^��k����x�xG���۵z ��gn�=4�4�	���WdM4@�肥�J�p�0u�xs�&q^�`
�c��><�$("�P��_��3�.�J�|�+��?�d���&��$ͯ���͂WL�!��{�|h���4�����M|�l~�1�:�Ω�>���U�_�4�0S�����x#�x���c=�ea�;y� ,b0V�u�Q��]7K�6�á�~O���-@t�/�W/S��8(�E���Kt㲬��MK�Lw¹��<d�Ji�];���w¹��<d�,��L��T^�`T�W�88�;矷p�]3t�}i�@�5�}�]������2���񥦢$'5�J�~���.����7�*���<�Hr��r�,z_�����9ƿ���=�Ҹ��tk@�Zۙ��A�>s��Y�&�������t���c����)��Y�6� ;h$	A�J�e�!�c�A�L'ӸT�?��i��N�N-��;���ݕ�
�o�`w����:ը⒍~����\�d1o�rs�i��5O
T������c�v�J��sr�l�k]m��2��+���O�ꢤ�Og�C9r%e�X�m��{��5�<} q�\E��0o@aT�\ө�M��%LS�I����5��d���zj5�Aɀ�� A�ST⃺��<kPj�^��3�D�I��
�[��b=��|�)՜�4�vIn���E��O�z�ώ ���]qI>�`��+h�5,Wlr�r%)cAQ17�b����#g�k��X�C���������C��֑xGV�[��WS�,�j:&AԢ�a\�DW��E��q�����C��֑xGV�eU���(�͊����ss2����`�|��K�z>���@]��8=��2��3�L����e�eV��iA'R�	.s�b��O���P�|T����E�E��3�L����e�eV�M�z$��P�^�6�V���l�p�H1�a-���7a
��r�S�B+����;��|B"�2�,.�Rg��L�*������5�m�bu�rI>�`��+h�5,Wlr�r%)cA��z>9�R�#g�k��X�C���������C��֑xGV�[��WS��񔖔�c�fi�d>G9���ļ���/���b�Bϱ��3R�e��ł)w���m�±��m|J�}�֖���J�_��e����7���{r��f���꜅�R��ӟ-�|qU?R�f��gn�=4�4�	���WdM4@ȗ��ƒ�˘��o���FO�W;D���P�<�F}���V6��Q��&i��N�Na����g�6���Q,|y�����Y���ǡ�C�a\Y���[C�W�v/��1h=��|Ŕ��lZR����,�ǰ���!�Ab�f�s�G�m�~]187A�SWۆay>��k\�����ܿ�(����5���ռ�j����)w�n��ukh�¦���@��8����S���� "5�]h�' L� U��֜��3�=���Q{�1�a-���7a
��r�b��j��<�I7��-5l*���T�I7��-5��5Z�����L��c⳯���Eu��oŹQI�~�џ0I� X�1� �����b@c{{��
J�~���.����7�*���<�Hr�`�_��QA3e��q���)��j)yc�n�.�_�t�H2v���Q�[��C���������a����"�$k��,�:�N�*�x���D)��g�%Y��̗0z�cULj� 1ɡ��&�@�}�-��w��k]m��>=!=�"���Mڷ�l��)��'���Xw�j�7���3R�e��Ӵ�"�6j��;٬sf.�B'=�:�,�y&�/S!��4_���QR�Xe����;���/�kI��Aġ��������[m��3R�e���V!8P�24%6� �7��)Q�XI��J�)��yf���x�M�g�������*[UxG��
�	?�<�a�/!O���������T5��t�\��ot[�W��Vg��{�����$�(��n� ׵����:�#T�a��p��x+6���Z��~����p7A�SW���)�aO�j��&����KS'�*p��0���!�|~�X��˓"��0��HXC/���eV�
��e,OL���t�b�hO�^+���\5؃a~y=�,����ێ_ϞB �'@v
@�1�Xׅ�LN��A|���]}����xT���b�c�r�{jFKL���:�G�h�� oj�VO����+���������᥼�5�/͆�꺖Z(��:�l�5�����xn�|������Y��#�¡�kU�%Rd�B���^��5��f�
�7�gŢ���ᣊ��f�T��nxq�� +@���))P�����X�C�HC�|��dq9%��9.7g�t���<���/�3��Ay&<y�;��|B����N���h_�zG6�o8:4�I���c�90��c��qq�KX��ik���`+iYb"Όd)��i?|	.�4��s��Z���.TE�g�������(ӈ��� �3�c`��0��₎���Ȝx�5W ��̫(>��o��X[�QB���X��WG ��i?|	.�4��s��Z���.Tv{��lw	����,Ǣ�Пe���;u�4�J��x(�i��/Rh�x#�L_�(D{ͬ�y��IX0F�M�^����'�֫��XA|>���)��뮗�w�ތ4�7�K�Š=ԕD��6c��wV��߬�F�<�t�W(@M�(fw���'�̗������k2m�;��|BG�a�����C1zh{A�dha#4��������o�^Һ�^E4+у��b�Bϱ��3R�e��ł)w���m�±��m|J�}�֖���J�_��e����7���{r���i���A�* ^��\�v'b�'=�(�ժ�E�$��*�]u*+l^�V
h��,��G���۵z ��gn�=4�4�	���WdM4@��&����˶�6�>��ʬ���7���{r���i���A�@[�_zβr��o��SO�W,�P &�\iT�������܏g��L�*����`w
��Օ��qvdЧ^{�jM|�"D^���\�}6��~p�=�J����6x�F�-LU����{����J�^��4br�����w�����P�<�F}���V6��Q��&i��N�N-��;��M�z$��P�^�6�V���l�p�H1�a-���7a
��r�$Dc~4�A)�V��/�����;٬sf.�#@�Q¢�r}l��L�e�+S��2v�C�|J3J��$5w����k��뗁��cA��짦���O�ʦ
���c�v�J��sr�l�k]m��+qO1U��#_"`��Rss2����`�|��K�z˦9��iժG�p�P��c� V��	��yv�ʯʗ�bu�r��c7�
W���ݤ�E��p��4#h���C�m�t�T�.�p�ݷ���1Kޑ�l��'�.ᬵy��̒�R�K!����� hbvk~�#xXX�dPh(??�d���&���xBS1Or}l��L�_�Źz=+��T����oGo�Z�������/�)��ɖ�c������+��?G����������!�2��~;-;*�7��vє�&�������7���{r��W�Ty��5��D5lR�^Ƒ���)ύ^��R�^Ƒ��YD�L��G[�� ��aP��k���[!��eC��[�����p��@LV�0L��{^{?	�c;@D�
��IouX8�������=�Ҹn1��Et�!z�t)P�a[)9b�jT�.���I�]�Bbr*N���)�[���6�5�9�(��H��Jy`�����e��+�ה6� ;h$	A�J�e�!�c�A�L'#.�YS�J���֑xGV�F�m���}'!��/������ٝ��AL����	'B�ɏ��]�!��	Ǹ�y85��^����d��;٬sf.�#@�Q¢�r}l��L�Kp]k�sE�z�'��4_���QR�Xe�������(2��&�;�*t5����J#Q��d�)bU����,Ǣ&n'o��WcUB�J�-/�)ع��7����]F�L4=�m<����6U(�<"�͊�����֐�f�-Tl���a[�{��+3?���*��+kt�Oz���,�ǰL�[��V�6�V(>�׀��6���pN �DؿZ���X����O\<��#���FQ�Q�I��o����De�A���ۖ\H|J0=�Q��Se����4�U��O?`�����R��󬽋?V�ҁGG�k$��"T�g�0�u���U�u!�?8��Cd[UUt�\����P�]��w]3k�ul�W����nF���<�W�.�P��c3���3M��	��3��a���!@�f")Ut�\�ASU�
T_�mS8<�n��._(������[m߁��(2���M������'�u�#�%��>�r�.�kRc�}���Fo|k�Lbx(�i��/RŻ�&ǥ�̫IX0F�M��D]�V۪	�}a?�d���&��@~�,r}l��L�/��*�H��	��e�YV�����a�:�?J��v�#��#Z�j|�>�O򏇱�{�� ,��rQJ�ڣ.�����2����v�x�;��c�}�CA�2��,�r�L�t��n',Mn�Va��G5����k:���"!9"X|]�c��%#�N�ǁ�f�T��p_U
#;��|B4���,����c�}�C��2�������t��P��M��%LS��b���jp���gL��P�����,�ǰ���l�{��4�1��3�MY}�!S���htam���M����A�m�(��D׉��h�#g�k����awf�#�%��>�h0Z�W��2N!�y{+��VӁa�|�4�b�6j�"Hsfw(��-O�#�58W�����,�ǰ�-M�bRr�a���hJ�����R�/c^ׯ)[�de!:�^�y�!B,�1�J���S�[Sf�;B�A��Ja�'6���L���Pe1��*����:ߕj�={"��s�-������X�m��{�6;���D8��2N!�y{+��0Ex���X (�M 0b/0�X�m��{�Y�l���^�v{��lw	����,ǢL�E��<U����;��|BF?U�&K��"�9��J�j_6A.r?!��W���r|W���/;��|B&��im5�S;�d�E�H���A^A�sO��U��-ȼ[�˹��K6"�%��(��v�r�i���]�C�;�׀�q�R�āy���Rkj}kqx�>yM�Ñ�j�v��"x8���¥��w��D����D�G#��Q������ssY�Kv�c��Q��"��0��C��-��K�E�sI�I))����A�m�(��nb��I5�4`UV#-�[ҭ�Ă~�*o)�Ylom;���'�u��1�+5����/O8���j|�>�O.]�H��~�1�W���&�K�VF�]X��˒�Û���G�'����w=G-���m����>Vu���d��sR�/o�)���)K��I��>z�Vg.N������[���(?�%WJo��_�n�To�[�C��-����?����X��kRCլ�=`/Q� a⣃_BB�"h��.W��z�h1Vc��!�^-I�!A(��&O�a��T�0cU;�^P�G�ℴ~WH6�	���N+��������T���<��wn��A'@����/�$z��
7�g��lU�h�Rv"4a�,�R����,��Ĩ���pZ����
�+��Jb6�3�I�M07E�_��Y�Rw2Լ���.��;L!�����k3H�)�.�-z[�#�Q�le(Ԁ�?�d4)�Ubۼ��n���I��}|k� 7��q��0�_w�b,&�N�j�a��I^���	0̧�LJ�C �\���ssY�KJ�	�LÆ�b���[Q���H�V�������[b�����V�I�e!��nH�W��ž��v��V�y%�ЧX�m��{�b���L�>j%J���E[z�taS��R�Xe����b�A��d8���������p���+cErR�����,�ǰ	M,��rER<�v!��$�a��{d�v��X��VB�����#���FQ�Q�I��?�d���&�8V<�V���A�\>W�/Z��B���[@;��|Bᜮo{Q��ȷ��>m��Iu�`�o����[m��3R�e��.]�H��J�ڣ.���=ev��=�֖�QБ����t��h�	�Ȟ���?{W¿pX;��|B�����z݃���,h���w*��	� ��z� ��wqMYxw��7�ํ���Lu���g��n%[��t�$�X_�x�������Е6��!�G�ݙ�Ih�	�;WE���?nh�5,Wlr�r%)cAQ17�b����#g�k����zb����2�ę�u'b�'=�(�hU�AG��iŞ�W�%3AԢ�a\��?�D�p&��2�ę�u'b�'=�(�o<4y���W/S��8(�E���Kt�m���i�s���1�R�n� �}DG�;֬������8=��2#�(�>^�l�'s{	�h�v1a{J�n�G�����P�|T����E�E#�(�>^�l�'s{	�hj$��1�#tss2����`�|��K�z�
��vK���p�+m*��"Ϩ+`�|��K�z��l��jV��	��y>��
6��Ih�	�;�c�9�,Mb�f�s�GWE���?nh�5,Wlr�r%)cA��z>9�R�#g�k����zb����2�ę�u'b�'=�(�hU�AG���i�<�~�yâq�t�d����x�K���P�|T����E�E#�(�>^�l��e�eV���W�O�힬���7���{r��f���꜅�R��ӟ-�Wڭ��h�Ɛo�c�?EcD�=1]M����_���|��
�|u='�c�-��;��F��zF�ۗ�
Rۙ�)S���%��V�c���cA��짦���O�ʦ
�[�s���_����J����
i���R|�1�a-���7a
��r�$Dc~4���V�ptj �0tw�*AI����ݴC`��b����^�;��|B������+�+\����[n���"'��l������O���FW�&k@C�Ɨ0z�cULj� 1�C��(3��7�q��J��v1a{J��)���H��ɲ�cz���ł)w���m�±��m|��������!���c�A�L'd[�L"[S�|u='�c�-��;��F��zF�ۗ=WEڠ�ܣ����k��GJ�v�m��+���J q�v����6��w�1�l�$y��t�iZ]XF�hx��G��S��Ǵ��BR�^Ƒ�Ӥx1j���k��!a�tc�&ck��Wڭ��h�Ɛo�c�?EcD�=1]%�o�.���]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��sI�$����G[�� ��aP��k�= ��j��C��[�����p��@LV�0L��{^{?	�c;@D�
��Io�p��76,�/^;؊��G���V�0L��{�*���<�Hr���Q,��Б�����Y�M���˻��0y��<L(\Ӧ�ݡs����̲�2�!�O��V�/�|u='�c�-��;���֤���n��/�����~�X����ɲ�cz���Ӵ�"�6j��;٬sf.�yWL�l)�q�\E��0�-��*�6[�j|�>�O�u�Q��o{k�h�+�d�)bU����,Ǣe8Υ���V4%6� �7��)Q�XI��N�#{Z��M�g�������*[UxG��
�	?�<�a�/!O�C�)1p;�V��ЏL-Zb��T�Q5:�?J��~AP��'�X�m��{�b���L�>j%J���E[�|c���r1�1�R���'p�iSq ^��y�C瑘�y�����[�/��2��_��෧0��ؗ.$!��C_Ec�r�5��]?�����e��eK,�(���B��D ��jA�48��U2������7,D{l4�~����0_�	k�JA)�v_���G�ԝ�K� �2�>E�p��m�Q� �l�V��Ys���Eyֱ�J�y�y��_&���y�	���Ԇ��΋��[ޠ+�����gr4%ܔ���	0���=ѿ�wf�C���	i$�s���[14��6�z����dI״�`�'�h�!�Q��q�D|�Q����[�/��2	k�JA)��5)��y6΃վ��E5��[�~2΍�/���ʲ׊��ֱ"?�d���&�w׶bZ"󞶿
�]�ٹ��d�
�4"�9 \�Ԟ-zq8/�
QA�y+��A4
�t�\��ot��v�02+߇�C�q�� w�wAk$�V�a�g2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!/��KJy����YVctW��X=t��w���'�G��49�V!��#%�/��Z>LW� ���bs_W7�]��m%�/��Z>L%C݇-�%;��|B/B�Â���&S�rD�1�:�Ω�յ�'�)���Ҷt�|��ޣC&t�iZ]XF�hx��G��!�`�(i3n!��i+�ť�n8���L��g�I��RhF��ղ�^=�
t�zg��p��I7��-5l*���T�I7��-5��5Z��·���~X�~���$^!�X;p`�����?�dv��oTN֢&@��&��|��p8=�[Ǵ��p���@Z�_F�k-�H��bf�?ǉ�=�|�)՜�4z�Gb��P�!�`�(i3|w�{P^K���3�<�p�� �&���ç�A!�`�(i3�\�!wn�ř�3�<�p�� �&f��vA<U�=PRpY.[?V��j�cZ)[���F	��7��z_nÑ2h�-]�o�Mt��1���(Gl�q�X癌��� 
~�F�踫g(�r�N�ǁ�f�T��p_U
#;��|B�w,�O�`{�3Vg���j�Txk^�� ���R�^Ƒ����"X��[ow_;O
�xkx U�_@�]t��fg��������B�â2N!�y{+��0Ex��L�.��e��~��������Tg#�o Yt��}��z�S�T�٥��T��?b�t���6����H�5�Y�w���bʺ��)o�N��*M|u�޽�vUM��)�� Ww��Il*~IP���*��N�ǁ�f�T��p_U
#��'8��)���"5�o٥�i��ݟ�^���\�}N�#;��=��ծ�+�� mv{��lw	����,ǢL�E��<U>Hp�y�7Dl�ggi�S��w_��Gb��VH�p�-a�D͢?�d���&�D���ƨ�w]r���nX�i֝�G\ibE�G!@)c�,���M�*��ud�H�A�m�(�����Y���h�ӵeo�;�iD�m;��|B���X/��əS\�R��)�POۭ�نL�t��ni��:$��28��p�!���V��	��y���˳���~�޳^���������G�Ȧj�rZ�0m�\�n�8�Z�Ѽ՗�zϋ�,n�8�Z�Ѽ���9$��H��u�d�ۋI7��-5r�p =(��8�B���ow_;O
�xkx U�_@�]t��f]���^��m���PH�F��׿]=ͅ�J<v�N*�9�c���kb>���pۀ��t�~x����J�u;��|B���0�2u��/n|���<Ӊ��S��A&Qne���J�";��%YM�ξ���I��RhF��j���W���?�d���&��4w�d��˩���.pՁ�=�nlTU�QY�O�5�%]���a(􆿳�k��q��־�E�&�y+�.��.f�Cz瀿3�_Ï_&-T�*�7`����M�Z���	s�����ه4�tZ�=��ծ�+�� m�ݾ-/�;��|Bnf��;�\sf0�s�I�c���;�z�����S��A&Qn�_��1J���t����M~V��	��yޮt
0�_����s�j2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc4�`�(H�Ps�q�6����4�G-rx��� 0v��W5���i7��0!�[�0>�
��`��<�
�d�ξ���Ix���Ka���\�Q�b�#g�k��Ps�q�6�f!��������raǹ}���,*r��`�*Ea;��|B���J����}ָ� ��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϱ�y�Zk��5/��33��*�	�ػ/W��^{Gj��J�1	�<����to��y�[��7%^�W+��W�
cʄѓB�@o��[ea�8���B����g��Tݭ�EB����1������L�,\ަ�It��+g[����=�-�o&l������ݥ�7�r�&U������G|M����6%�a|�\m���j��&����i�\�{q����W�Ty��5!�`�(i3���gRI/b�]6��e,fi�U�ž�'�t_���NDa�zg��p��I7��-5Sk��?L}Vx�%L�I��J)#�Z��@��)�[���6SN[�ZǪ����}�Z�!����2�R��!(`濸!�`�(i3Ĉ���rl�����@�u��oŹQ2Y��kک����Q��K5���Adu�Bg&��C��[�Do�9�ݚ�Н�8j��zJ�U<�i��W{���铸tC�8�J�Q����q����k��,�:�N�*�x١w��zj�R̶����N�i����b�'Be����s:��i��NU�q�\E��0	ozqP.!ū�ez�,�۞��	�|$�kJ��_F�k-�H��bf�?ǉ�=̇i�d�?��˺�Q���f�?ǉ�=�|�)՜�4�vIn���Q@w�w�SB}j��)~�2��J�J��
UU7$^tjn�jX���Z2el�ߍ���y�C���C�� ��@2�7�Ap�dp���t�u���-���c�qDrU��*W�q_҂T�q�w���r�&U������G|M�����ڀS��d���!iշ���������j�Txk^����2��'B{q����'6���;8=D�P�E6�k��q��־�W+��W�W����G�iA'R�	O��cb>��POۭ���Ɔ �����Vd��0�| ��HN��R��?�d���&��|��Li)����	C��F%�X��+M�ᴰ`��Z�^����	�hS3y�����ϲ��Vo[���˚����Z�ם�.J7h���/5U��nFW�JyS�N�*J�X�$����q(	�fw�R���ykb>���p����9�d���V��	��yG��Γf�-���c�q����Ν(�JZ�Vk�;��|BMR��P.��=�Da�;)�bx�Ω����
T+Fb%��C��:O�����z���AZ���d���!i�\>�ʘkN�]��0g�~��X��r:�G�?�d���&�`�Ӡž.m1)2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���B��I.¤�l���R���V����������q�©��'w��
�fʖG�œ����s��3�mAR�o	%�ϸ��#|S������3[�u8���иܖ��Q�P���O��a�����(��ԋT���i�@�>�i�ۑ ��� ����H�ʱˡ@^�N2t���M����V�܄WD��|���,���9^-�Q١Ӿ�$������i��X;p`��w�f���w¹��<d���<
DN��X;p`�ct�:��RE�QS����>f�?ǉ�=Vx�%L��]n���@�����T�v��1���5Z�������/�U��֜��3�&8�,��ܠ'h|��W�Ty��5���}A�:�ߘ�)�I��<
DN�xj����R���it	�TU����z~���MK�Ls 3�:��)�[���6�&8�,�¿DĢ�WZ���q�������ȍry��	Gظ0�����@;w�$C,0�?����_F�k-��&8�,��Q�L�������!�`�(i3z�Gb��P��2��}�������Ə:S�.?<�:�,���P�,'"�i��NU�W����GS�*;qܫN�i������"� ^ŭ��S����3]]ҥ)J������}0x��� �?��$�/T�{0��d#�g�w0��䎀������p�2��}���/�^��-�����*��$�q�ʋ�x�h�k�t]�<Lz�l#�V��H��<�C�Ar��� f�Nd+l��p��;z�_��s�֙R���Bk�d*e��\@8GS��`n������ct�:��RE�QS����>�wo��Z��Ac<�p{�5�O�%E#P�P����9��g�ܧ*y*J�X�$����aV}�������,���1����,H/������,�ǰ�������'����2�,bxqX��g�9��,Y�����9C�������u8q��ǵc��5�%]����8�B���ow_;O
�J��:���闺����ő��"�\�!�{~����DKY�����|f���+X�E�k?�i2�.[W�w��fD�g�9��,Y��(c$�,w�R���y���,!��HC�d��g7,��(&���X�Ɨ��[�k�l4���Z_c�����o�.�����`pe�1	ٟ�,+$\�M�����p%\2�T>⺾�D@s�i�	����J������Ҭ�0��k��԰�/"��nH�W��ł-���������.��4�F1���g;��wT詊�H�V��=�WK=ZȂ"v�(=?�w-��U��)���Y;e�iKI/B޾PԐ#��go`iI9�o��|#HK��A(�c���_G��Hb� h�ҩ�!q��V��������ߊx#Q<Ne��0�U+�qbp@�՝� s�#04~B3��������h��`�����y_�mS8<�n���F�P�7��S��h��d\�����l��=�O�-v�*_�mS8<�n�ݚ�Н�!q��V��������:7L����(����C>:���[P�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�� �ѕC?">}���� ����!�@[�_zβrE��g�HbDR���6=+ڇ\�(& �����e����9�eF����k��԰�/"��nH�W�v�7�� I�����.��4�F1�筸b������H�V����GxE���8�ƌF�8;޶��*�\Q��,t�t@[�_zβrE��g�HbDR���6�ܼL�� iI.s�j���3�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ɸ,ǻ�|]η���7�,��n6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3��?�9ظ��ʱ�_ryhg�t�s�o�b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���a�<d�����r4���'k�����I0���ԏ�.fOe	� 	���R�	ڹr����hi�aDU�G�a�E�}q^J=����x�ԉ�>T۳�͕���׵���G��[�f��
������q9+t�}�P�HS|�O�D mWN!�`�(i3��?�9ظ��ʱ�_ryh/������V�>ȿ��'�8�nb �z�g��U-�ew���7Va��G��5���?�1%��?�9ظ��ʱ�_ryh�����˨g��U-�e�,���6+�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�T�t��5������$=}ݷe[u�;0��`��.��G��[�f�x���w�b��G��58��Տ*=��S�����u��Hic�{0��d#�����:%e����1�:�Ω��x[,�Ns��{0��d#����q6Ŏزm7Z��'HY-��^���!�U��}�o���#��Ӝᘡ����S���� "5�]W���`moF˯�+)��h�\ƙk����p�><��d5�:�w�+���LQ�/��V#��-��V�/�Eԣ5��)��j�3��	t���٫����'���$���k	�� L$g�(�Օ��qvdЧ^{�jp���,��H����8�� ���dp]g,H����N#=i-��z;���!��@��V�/�kt�����P�i2s��Y�7#�xIvє�&���Q�%�+2�j;��q,#�,D�t�uZ�v|�eY�6WffC` ��\U9����u(�G�&������ȍry��	Gظ0�����X;p`�l.�	�C�3Lv	̅��!�`�(i3>N0Θ��;b�-�2�>c��?Ӣ�c�����~�W{*T�i�������y�7/�YI#���2�:���f���g�4������S�|J�X;p`�]���!E�r &
�$Jf�?ǉ�=\.�l����k��r�a�^��D�i�ь�V%�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�*���j��jR�o+ͦ��t������ׄ�:�CTt �\ ��q<qs�B�ӵǶ�	��l�N[�-e	�z�2������A��<��T0���S=�Z���6h�����s��Q��sr �����c���#R|��\�ݔړ��0������Ѿ��/@�Yx�զ��eY�5��R3х���W���Bm�����y�3t�ʨ�u�w�@��\����*-�,���O�]�m�w���i���Z����Q�Y���*��d(c2g]=�v��&x�bq+��T����~��@�.��#=b|��ޣC&t�iZ]XF�hx��G��!�`�(i3�(}y��������i�?d��A ��+���LQ�f�?ǉ�=G&%	��ڏ�<
DN��І��%n3������0�O���]�|��T�5�d�,W�hQ�GvE��?��%��h�r�|6�gb��A�h��+FeA'�u���}| �e����kn4@Q�/�!�`�(i3k/�z�xEQ���*[UxG!�`�(i3���ꀍ�˺�Q���f�?ǉ�=��9��稕C��S�w��iY�;����2��}��CϾH�)�h��=;�)�^�\q�\E��0ס�Wd�#jsrCm�k��/z*x�n;��|B_�&F���b?,s�ca�$G1�O�P�9�L�,���F@;��7,������Z�׽�刍X��!���ū���t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��0���ɥ�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS�)���܇�a��o��ё\Bk�	�Ni�{�����f[*b~*��s��,l����M?��y�!�`�(i32W���R0(|v��t�a�^��D���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M|]η��q��_N�����,�ǰTm�v��G�g�v��Z�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�Z�@ns䟳��LQ�%�+2��k��kK�I�Q4p�/Cj���C�1,�A��#�jV�{+��i�Iu�5�O�%E#P_TR�\+�[�ƪe�0cwU�R?�[6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3e�v��ҵl�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS��%�����d��-��![L��^C�+a��o���H�RtV�^�3��C���H�� �YߥթD�[*�Bi�v�V��'�njVfV:)��{D~�u��r��!�`�(i3e�v��ҵl+��%�k<.�B�0���;�¬pX��g��U-�e�,���6+����%>�rGO�D mWN!�`�(i3�v�Wס���G�K$x/��&���Xd	�/I%L�Q��T��� h�ҩΪ���l�� m.x��(��p���'jsrCm�k�J��6�d�C�
���W��3��ݪ��=��l�r|{�,��5�Q�J��6�d�.�B�0���;�¬pX��u]9�#�I�s)l໶�,!�`�(i3�W�7�tM���p���'jsrCm�k�J��6�d�C�
���W��3��ݪ��=��l�r|{��\��~U�J��6�d�.�B�0���;�¬pX�出����mo�B� �b��!�`�(i3?V��j�c�:#��XB��4,�Q��U����z~��6��	���`y����ݚ�Н��Ra])n#���r����!�`�(i3:8�zH_ɗ�;2V-W��	c@�^ k�1{&��� M?��y�!�`�(i3!�`�(i3e�v��ҵl�]�!��	Ǹ�y85����[��xԲ ._�U6�bL�f�z�����jV�{+�fbmDF�!�`�(i3՝� s�#���k$ !�`�(i3{k�h�+&k@C�Ɨ0z�cULE��K3�j�U�V������:��`6;�¬pX���O��R�^Ƒ�ӆ�v�9��!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j���_J��`U�a�(��^GѬ�_aT��3G?�d���&�����t���B8궩�t&%�=:���'��-�3��#?1�U���gFck
����ɣ�<�f��jV�{+��i�Iu�5�O�%E#P_TR�\+�[8$u�Ӵ-����t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��04>^!b!4b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3��Nh�=f[���������<�.�����8��GM��-����!�`�(i3e�v��ҵl�]�!��	Ǹ�y85��r��3��kO��u�+�uB;y�cU�^.����P�7� �:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�8���SY�N�xʫ�A���;_��8W�w��fD)��J(�92�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�D� �B���9�V��r"nq���z���;�Ӏ�K��tV�:V%�&)�򄭩I4��欱���j�����|��ȤDL�>5�C����A��,��I4��欱���j�����s�QN���d���!it�td���52�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pdl2����}*X�K{�(��	}�@�r�<Uee�N�����0�=��;��|B���r�����z� 3P���@{2귑����Sa�!�`�(i3!�`�(i3���i����k]m����}Dq�f��z� 3P���@{2귑����|�kI��RhF��U>V%`�~�߇���t�k]m���E�i�m}66j�"Hs�@��C�,ԭ}3Y�Z��E��3?�d���&�Û=�������fo��ZpW4%"������k�I��RhF�䦓����������A2wKaC�IX0F�MV�ҁGG��Ւ��n�0 zK<U|r���3f�\�J��ײjw�ME�po守�ubs��2[�a��o���H�RtV�^����lr�{��|e��0�U+�qbp@���\ Nhk+Q�h'�Ȝx�5W ��̫(� h�ҩ���fCI��8��GM��-����<�6�Q=�I��� g~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D�Ϛ�-����!�`�(i3�Y�
 �vc�jj&��G�9m6�̟�1��"~6���aq��3=]��m�D��-����!�`�(i3-3!E!����Bf���̓@?5ɔ��,Vr!�`�(i3��Id�!�`�(i3�XW�����5=��)Q���nF���<�W�.�P�	��
�Q�}<�6�Q=���F��O��ݚ�Н�烉s)�v�bP�63Z�t��Qѳ$G��A0ok��烉s)�v�T����� Ԕ׹�ն'�U;|�� �Rɮ�/���¨}�n/�J����lh�o��_�Rv�䩲$��ƣ�Ę�2{y����i�q,?5q�+�#4��F��8M�po守�ubs��2[�a��o���H�RtV�^��KV�9�]Kߩ�d��my$�N��o�/���;�I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^���9���LQ�/81tSjv��� л��"�Nm>Ǖ��U�._�3
�v�v-}�	mp
���U{���8^��hJL��;���N�4��N	�7q������O�޳!?�R��n}�����H�X��WG ���N��b���c]p�5�	$o��Z�_�n�To�[�}�~��lg�7&�oe�XƤ5_���M���R��ӟ-���J��RQH�RtV�^�XW�����ZRR���dN�<@Iv��nt=:��:5A��p�I��Yq���k$ �� л��P�궊�2�����8!��?V�&�2���)x�?{���x.�Knq��5+*��4br������Ľ����Չxv��Օ��qvdЧ^{�j����'�����Z>ؼ��XyH�RtV�^<�6�Q=닓.�`�33c=��u<Rleށ�!�`�(i3��Qѳ$G��A0ok�®� л��5ߧE4��<�6�Q=���F��O�C#/<���q�5ߧE4���Qѳ$G�φ��<�6�닓.�`�3����΅�yǐ:�̋�:.�{��T����.������胋�M��a�-V�Cp	��?�?"���і�O:찹��S>���P��Y1C8�L�-�zm�2����~8GJ8���,�I}�F�y�^	#�-w˕���k�S���ld �jX��b�����ݻ��"~6���aq������J�?�d���&��������꓂O�q��.�1�4�o� c ��*�O.�N��A$�P������5d�������)G�9�=�1��*�
�I(͂X��WG ������&�Ko���&�@�}7�q��J��v1a{J�h�µj�!{�N<'��Il��!yZ�d/�����C�V���3��ֳ�Ե�i ӫ/��mR�MP��G�>��jj��r����.�aq���XF;�p)��
ۼ���Xv�"�M�)u��)o�0�ʂ�j�Ï��	�l�lM�3 �\Bk�	y�}�6f&r#o�]�ʄ�q������O�޳!?�R��n}�����H�X��WG ���?�,t�J�}D՛��W;���\�H��/Sg�w��'o�MdGN�������m��8\�Ia#i��N�Na����g�6���Q,|��,�ϣ퉧:��oQ�|i��N�Na����g�6���Q,|h���fn�g��]�J*�Rs�08�b(�����̜�I0���ԏ�.fOe	�HlU�!=���~�����gn�=4�4�	���WdM4@�肥�J����V��)x�?{���x.�KnqH�Ћ�r��%�z�J��z[�A���3�L����e�eV�M�z$��P�!�A˪[	��j"jȩ�i��N�Na����g�6���Q,|h���fn�g��]�J*�Rs�08�b(��R����� ӫ/��mt���������m���šB)��zR���b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$A�׭�%*b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�/%\��jX�m ޶&�hbvk~�#x�%��4�w����m�����F��O�n���šB)�X[��:~6q���w�=��u���'b�'=�(J�}�֖��-�X]t$IDW��E��q��u���'b�'=�(J�}�֖�
�c���zU���̜�I0���ԏ�.fOe	�HlU�!=���~�����gn�=4�4�	���WdM4@�肥�J�h@I �y ӫ/��mR�MP��GX��WG ���zR���b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�V�һ�d�#P�j2E�?��Id��o<Z�L5a�"Pn��s�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a��Mg.6�k���'���o|k�Lb���'���o|k�Lb����k��?�,t�JN��	�Ȓ�cЉ�M�K���]��i�a�sir��5��܊K�+���w�PjI^�UI0���ԏ�.fOe	��<������r���3�:�����{~㽕���䕽v1a{J��=t�z/�����C�V���3�O��+�El�n�.��ɠ4�04�jf�nٚ�2�,�n�.��ɠ4�04�jfc¦�.��aY8.���׹��*P�{��	�ɭ��
/��y;��=�m�W��n4p�`6j�"Hs��Z�W����/��hH�C�F?�������L�����%C1��,2�A���ۖ��S�<Ԣ�,
�u#���n=�Z��W/��WuB=�r����'����IX0F�MV�ҁGG��ABk@�0h�5eצ'ž1�|�'����Ut�\��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�V�һ�d�f��xp�M�C�x!�H�k��^)ҠN�2$�I))����A�m�(�}gQp�3+�\�G�����dc�@c�����hX��WG ���͹�k�9��d��-��!�L�F.	-�L��&PY~�y����o)�T*�c��܍w�S}�u��XC���}D՛��W;���\�H��/Sg�w��'o�MdGN����9�d�L�c]p�5�	$o��Z�_�n�To�[�}�~��l c�o�u��.ᬵy��o"#}aUt�\������-�G�h��\`�R�kA7��V ��݇!�
D���;�g��ޙVb�"�I���I�����OeU���(;�~1��_���̙�R��I���I�����OeU���(�&�r^-���.������v�8:������fI��jÇ+�_�n�To�[���9�P�4vE7�MW�o�>>����I���I�����OeU���(�G%i��A!��: ��ao.\C�kG��R�	J_g()��ikp���H���F��kt'n
V~$����4~V��3�L����e�eV�M�z$��P�!�A˪[	��j"jȩ�i��N�Na����g�6���Q,|h���fn��0h���J*�Rs�08�b(��un��7� ӫ/��mt������q�)]Q�x��r_��mzf	�$NT�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a���4�M1��A���ۖ�k�V\�#P�j2E�?�5ߧE4��>je`��@d:�����{~�Vb�"�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a��:��O�?�I))����A�m�(��C��AF�Р=��'e����&�@�}7�q��J��v1a{J�h�µj�!���5��Dao.\C�k]�	,��QUt�\�u��a��i��N�Na����g�6���Q,|��,�ϣ��19TH���"L?�����G�\�4���gn�=4�4�	���WdM4@�肥�J��eqm����gn�=4�4�	���WdM4@�肥�J�:�D5��h7�xȀ��D׏�����Mp�-a�D͢q��`�L�5ߧE4��; T�����8��GM�v�]��1VTҝD!u�Z����pG�p�P�m��������a-6�Da�K:+>N��	�Ȓ�cЉ�M�K���]�����` ��y/�����C�V���3��ֳ�Ե�i ӫ/��mR�MP��G���:��KY�[b%Ɨ����7�P�K�+���w���řA{���C�x!�H����'^_J���|{�mdJ�1���)�@����p�-a�D͢fU�9�׏�����MFi��|F�}�WP']��6�~����0D�N( Q���L}��M�~�ajJɫ �~wS �X�C���������C��֑xGV�eU���(;)(F�T�	�_��:��u���'b�'=�(J�}�֖�ت2�<�O��gn�=4�D-'��7�q����r� F�3N�����	��gn�=4�4�	���WdM4@��&����˶�ּX�b��c�fi�d\'�s�@#F e8�~����t9N\ا��=tu�㺅ڐK���l_��`N�z��7|^���~�@3�$��I)p�z!��U	�`�o��_�Rv�䩲$��8��I��.��|ȃ�A(�c���_G��Hb�wd�#<����Tk�-������c�����B)|DՃ���lf^�;��C+�G~���M��Nv�*~A�,��`������]kK�+���w� �s		��N���u��v1a{J�@<}��A@g()��ikp���H���4�:s� �q��]���~��-Y[;�wQ���սv1a{J��z*  x�I))����A�m�(���}܁'�O��<��J*�Rs�08�b(��l`��\1S�u{hK�'��݉�=�����w�=��u���'b�'=�(J�}�֖��-�X]t$I$�D���O�J*�Rs�08�b(��p�QD�á��&�@�}7�q��J��v1a{J�}D7B��#��M��hbD��ڙ�n�ZLN�	���}���x�A���ۖ��1�:��^ K=�b��ġ��,��{�	���v�8:?�'���&!����-�g()��ikp���H���G6.�~�݊���w�=�����C��֑xGV�eU���(;)(F�T�@Z
��#���Fi�"τ�����p��}��aq����(
}���û��i��N�N-��;��M�z$��PКą���g�U4���Z�Ϥ�h��K�r�\E�6O:��2bv!nU��K.��QW�4��i�P�
ɴ��z�4�	���WdM4@���d5���J*�Rs�08�b(��R����� ӫ/��m� ����+��J>�߯�"5�o٥眣TFC�)x�?{���x.�Knq��п��Tg()��ikp���H���G6.�~�݊��n����,6��œ�'�����Rkj}kq�MT�5�o[�a��[�s���J��sr�l�k]m��8����`�'J*�Rs�08�b(��R����� ӫ/��m� ����+��J>�߯�"5�o٥����Y�JM�b��v݋N�����7u7҃Q*�6������1�R+-h]�83NI�����w/,g{Y#0����l��=5; �e�W|��6�C��(3��7�q��J������-VL�Q�K��x�A���ۖ��S�<Ԣ�ɨ]^(���Ѹ���_�j�`���: ��ao.\C�k���uf|ò���
��_������B�K��1��n�da�ۣqM��X�~ ӫ/��m�D�K����g1�#�(�>^�l��e�eV�>�3�eZ~�f�R�&Aju�j[����#��47�
ɴ��z�D-'��7�q�����*8���������@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*�Va�ir�4br���qP�V>t'�̗����S]�_�_��Ut�\��"�Nm>�DQrv����)�x�.���;���8$_Z
��9�#���F�H۷`n
V~$ą�m[���'���c�e�+���4.�*�l��=5;�a���8n
V~$� ����%��>M���b��v݋N�����ה��#m��`$�\�����ZLN�	���nE�g%�zR���bJ�%Ph�r^m"�OB7A�SW�N����4�P��/ ں4��VJΣ8��3�L����e�eV�M�z$��P�!�A˪[	��*3)�����3�L����e�eV�M�z$��P�!�A˪[	�2��h�d�)x�?{���x.�Knq��!cI͸I))����A�m�(��C��AF�Р=��'e����&�@�}7�q��J��v1a{J�}D7B��#��T��n ^��A���ۖ"'��&އp��;�{����G�\�4���gn�=4�4�	���WdM4@��&����˶O@�s��M���c�v�J��sr�l�k]m��n���=�y���5Lwn�3
�v�v-}�	mp��"����I0���ԏ�.fOe	�HlU�!=T۳�͕��~K
eڟ7���&�@�}7�q��J��v1a{J�}D7B��#��.M�LYq^���&�@�}7�q��J��v1a{J�}D7B��#�w���{,�:g()��ikp���H���y���@�Krw�&�z<a�4�ڈt�[b%Ɨ���û��i��N�Na����g�6���Q,|]���#��:��oQ�|i��N�Na����g�6���Q,|6.o�7�OY����A�b��v݋N�����|�+��)�Р=��'e����&�@�}7�q��J��v1a{J�}D7B��#����5��Dao.\C�k]�	,��QUt�\�zf	�$NT�I���I�����OeU���(;�~1��_��pPo��zT۳�͕������4~V��3�L����e�eV�M�z$��PКą���gƜ*3)�����3�L����e�eV�M�z$��PКą���gơ��^��Mrw�&�z<a�4�ڈt׏�����MJ�1����z%�ژ�(�*4��%�#o�]�ʄ�q�����Q%I4��뇿D!�0�?�R��n}�����H�X��WG ��W|��6�C��(3��7�q��J������-VL�*3)����#�(�>^�l��e�eV��_�vԡ3�OY����Ag{Y#0����l��=5;N�����O������Mc�WT�D�3����K�F��_�M8O؏����:�~�1ߩ���ZAL�:������`4��D-~nҙ��ș5*�M��1�y�I��m�n����[�s���J��sr�l�k]m���������N��-���'�[�s���J��sr�l�k]m��M�s�Ӟ*��"xC��-�T(u	M^)FU9����8BW�R7���r_��m��zb����2�ę�u'b�'=�(��$��O
ɴ��z�4�	���WdM4@�p�r5A��J�1�����u���"6ɲ�cz���Ӵ�"�6j��;٬sf.���Y�m��
ɴ��z�4�	���WdM4@�݆M�g���󑟇���-hbvk~�#x}���y�Db��E(�\�H��/Sg�w��'o���u���"6����׾dC�ڃ�P �J�bMfo{��M�M������W&Z)�8�i{2!�Mn�g�L�2w�f��8/���u"MP�UUc�WT�D�3����K�F��^VE����t]���|���N(�1[�G���Kn��ɲ�cz���Ӵ�"�6j��;٬sf.���Y�m��
ɴ��z�D-'��7�q�������Q�$Gu�w��Ds��>���R�^J|WQ	��2�b��v݋N�����|�+��)�Р=��'e�C��(3���-��w��k]m��8Sg��
Ԧ�C��u����1m�Ut�\�8�%<}���"'��l������O05 S�s�lɲ�cz���ł)w���m�±��m|�b��Č�?��|��袔MUt��!�J��Y��̵�"xC��-�T(u	M^��|A�I���pP�$D\��z�
ɴ��z�4�	���WdM4@�E�RN�- \C��(3���-��w��k]m��������C��uu8I#M{c�}���Fo|k�Lbx(�i��/R�;b�-�2�׏�����M�[�S�n�H�,l�����(4G��>�S���%��V�c��ݕZ����pG�p�P�m�������3�� �f������.S��X��덎a-6�Da��J6����"'��l����C1zhi�Y
�,�LٗH�1�"'��l����C1zhZVv ?JZ��,H���F�]	
~ao.\C�k�Y�\�n����[�s���_����J������ݱ�JGy�ˆn����N��+�CAƨ�D5���a-6�Da��zb��B�>��֑xGV�05 S�s�l�1Qa����˓#�������\|u='�c�-��;��>�3�eZ~����z
��|u='�c�-��;��b'�Y@%^~>��mJ�1���K���L���4�04�jfx(�i��/R}�	76�&�� Ӗ�t$�)�vxv���}�_�� �R�"�n)�Q��ܾ7�'��ܷh������{ԕ����D#8`�k]m��v��z_����6��Ɔ ���Ve��˅�:�}��E5��OP�Յ������ꏶ�Ij�'��щĽ��1{�K�f(&�/� s�Y�����0�;�s�$�������E2��W䁱3�}$}��î�Zq�������L`G�v�~��]X���k���_��&7��N:��"^���H> �([�4����tm+�E^J*�Rs�08�b(������T���n��<��%m�Y$� 1���!��|�+4K-��4~H�<�&��x����<�S���c�&����:)x�?{���x.�Knq��5+*�����˱f�렾����o0hp�J$!@S�@��NXA��� �h��N�Mܲ���C�>5�,}9P!��|����GuDc%^oe�Y��k���_��&7��^�F��vh^���H> �s�bͦ-(�Ⱥ�kJ��*���[�\#���Ƹ��p��6�>������n�O��Ե�Z+���g��o����>�/�d�@���G3��X&+M?�n��<��%m�Y$� 1Z�����j�r]��=�찺pl�E(��6�� ~^N�gG`	Plh�P	���Mcyö��]f�,"y���L? ���U�d�@���GU����N�="��u���܁�i��:ژ�����Z4GL�}�痽�����)�aO��������J�)��Z+���g��o����>�/�d�@���G�%�4�'S!��#����В�S���GuDc%^oe�Y��k���_��&7��^�F��vh^���H> �ݎ' w%g��_���cشŀ��`�z���xl%����v缐%�/�<�|K7�&^v� E#�F2~��E,};�^�)׶9�H*.埲���G4��cf�l6�L� *���˿O�F�{�e4���ҏ�n�%$3��)�M8��	��?�'��/2RIh���o��G9�}Q*%΢Ӟe�H5��M���*�f;!+�+$�����^/e��d]� ���_�hbvk~�#x��q��ZVT�x�"��XƤ5_�J�	�LÆ���#��}���![<"XC}ץE�$��Ly����:�����U��2�ڥ����Ⱦ|����?��eߍ��鋎Z O\������U�._�nQ�rV��q�t7�.��/��SB�/���\VO�l� mr�m� Z�l�o����>�/�d�@���G�X���.��ġ��,l5R?}�b�+��z���&�2���)x�?{���x.�Knq���'
�?��p��6�>z8^�G8Lu�>�� 6�o8:4�I���c�90��c��qq:Fa�7���W"�P�K��q��[@��'ž1�|�'�������H��e��k�J��ֽ�\����g��U-�e>� {�}���my$�N���Uە��jz�\=�/��8y����Y)�'�m���[�4�f,�{_8�Y��=�}�Vݨ��\9�oA�d��JXl'�T��~��Uг�|<������M���LQ�/8n
V~$�+�$�i4�ǖ��`Y��}�O���硙�t�\������n�O��Ե�a(􆿳�e�&���6�+�$�i4�� N٣��}�O���硙�t�\��������J�)��a(􆿳�e�&���6�5ߧE4��J�1���k_���b_���~�L*f3�~�;kΗ�31���鸗r�!��=cv6�Ɛg)x�D�����X�X� U�X���#g�k����?��j:���'�Ȳ��A$�P������5d�B� ��~��U��B��-ն'�U;|=�9U'��A(�c���_G��Hb=��"�ԭ��\VO��1��0����,?}�a�,��Sq'�@8�Qq���z���nF���<�W�.�P��c3��4br�����w������n�5�����}�pIɽ�Jz_�b_X�XV�b�z'hۉ)K7͍���E@�����s��U;4���^a�nu4Bޗ��jw�	����/�ciJ��Yu�����Fodً]�N� &p�ۻ�F'i0QW��8�	3i�\��׹��t�M��|S�/���[�4�f,.�q����e8�b,Qk^|�ˮ���$:N�t%��zxa(􆿳�e�&���6A�іx���\&<���٘ۼ�%6Y�G�˱�ߓC娤l��
�~�qYUS���%��(ݒ�hU�y�搲)���$:N�t%��zxMg.6�k�5ߧE4��rw�&�z<a��N� φ��<�6��PT�!�wd�1�D�V��	��y����U����鸗r?1��j�=�*%΢Ӟe�a�f+(��R}��ک��\VO�l� mr�m�(�s׷�~O���M3X/��A���-�Vb� ���������J�)��a(􆿳������>�,r�/<]mz�(�����2a� `�ئ��# ��6U(�<"��q�
�`�N�9�;�S��2a� �6�_��f�D�!$9�:�A��� �c�eC(�5_��&7��Ј-�S��f~��DV��O8Ľ-�X]t$I��6U(�<"f6�8Nn.�!�6UVo��6U(�<";�~1��_�u�9j7Zj�� N٣���RUt�E��6U(�<"�; Me~��?���J��J�)����ʨ )o�or�K��:8���+����d�]�����0\)����+�ڔ�I�����t�a,�$a���h�4h;D8���:���`�����O�Y�a�G�'������E�n���
Ո�C�hk��Y��A�m�(�,"��h�2
��F�l��=5;z��˻N�dLd�r:ha3B��*w���6b��ʏ��Z��4`��O::��n[I?��8y����i��?}�˼�f���MWdWV��	��y��I�A���U2�h=c��_���	���%�� U2�h=c���9�Y��v�c��Q��"��0��C��-���R��)�xQ�b��v݋N������Q���u��N�"9���b�=�`~G��?.�#g�k��֓&Zf��%j_H�ˉ���0����f�Nd+l�Yҽ֗�x�\c�5#�y�mDƝ��0vdL�_E�������,�ǰ	M,��rER)�H[ɳv��X�x�LV(<���wj-�::��n[I?����$ڑ�N�(]n�5+�D�k�x<C��:�c-yi"�����2�^˧��t]����ض?l�� *%΢Ӟe�a�f+(����&�K�VF0��<�@QQO�W;D�gL4�e�d�Jw��3�	[ZZ��-�`��W��D5�|��7�OT�,���q5�n-�@�4ڧ�<�j�k�����Z���%�d��:
�r" ���]'\gWg��	�Z�kfc�L�C���e��S�J\7!c�2�����U��\ڦ'ž1�|�'����Ut�\��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�nR��ړC娤l����pQ�q��!W�{_8�Y����X���������4~V��3�L����e�eV�M�z$��PЄ� *��eR��n�J>|�
#�`�^{��u�oDb_X�XV�b�z'hۉ)Ժ=���]��4br��L��_��R��n�J>|�
#�`�^{��u�oDb_X�XV�b�z'hۉ)K7͍���E@�����s��U;4���^a�nu4Bޗ��jw�	��#.w^�oG��8��GM/f��Z�~K
eڟ7���&�@�}7�q��J��v1a{J��(O T'Q`���$���^��y6�T���1���A%�@* ����c�v�J��sr�l�k]m��^~W���\'P�����M@�qX�Uu�T��3���W
�����4~V��3�L����e�eV�M�z$��PЄ� *��eR��n�J>|�
#�`�^{��u�oD�g�)�I�졉�&�@�}7�q��J��v1a{J�9�+J!��Q`���$���^��y6�T���1�����@�g����Ǵ=O�W;D�1X�iRd��D�����X���*"��Zʊӽ�����4br���v���R��n�J>|�
#�`�^{��u�oDE���7t�x(�i��/RŻ�&ǥ��a���F߸��S�Ȍ�w��ڷ�"�l�7%�]X����Ǵݵ��O��M`(繉�i�O��M`Օ���4���M���o�G�m�?���bq��;��|B���l
����>Ź9f���D5�|��7�OT�,	3i�\��׹��t�uDh/P^s[xkx U�_@�M��8S.�U��)���Y;e�iK ����)c���[�����3fEa�F��x�ޝE��A(�c���_G��Hb��a-6�Da�Ɔ ���/r�G�vH��~�.G�`��ٞ�R̕q������鷂�nF���W�_te*�"��?�.>#�����c�v�_����J����肥�Jӳ��n�5�����}�pIɽ�Jz_�b_X�XV�b�z'hۉ)Ժ=���]�X�C���������C��֑xGV�eU���(�˃��'�	3i�\��׹��t˔R��}K7͍���\C�
<r�8����H�v�ov�*�Y�G�˱�ߓC娤l��(Q6D���硙�t�\K7͍��|��W&":nv�q����� N٣�SG㴊�?����q5�n�JrPQV��dh_��tCdN�<@Iv��nt=:ྵp�!���k+Q�h'�Ȝx�5W ��̫(��a-6�Dae<�Ia��l�9W�a��=2oΠ�5�Y� u/2v:�v�H|���}�pIɽ�Jz_ꛨg��U-�eQ��,��ǖ��`Y�SG㴊�?����q5�n��dq�8���/�#P�j2E�?��6U(�<"e��w^9u�R̕q���s���4���܂%j_H�ˉE���Z�Y�G�˱�ߓC娤l��°������R�wX��)C8�o���C�x!�H��Tp�����5���7�~���=���q5�n�>.U$�o�N��	�Ȓ�cЉ�MMe9���ݱy�搲)���$:N�t%��zxMg.6�kzf	�$NT�I���I���C1zh�6���Q,|�b��暴�~���=���q5�n�>.U$�o��	�_��:�����C��֑xGV�eU���( �H^䁭	3i�\��׹��t�{ƨ��;N��-���'���c�v�_����J�����&����˶���n�5�����}�pIɽ�Jz_ꛀg�)�I�졉�&�@�}�-��w��k]m��n���=�y�y�搲)���$:N�t%��zxMg.6�kx(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}�|&�xVgY��m������L}�E�6�����>Ź9f�Ps_*�GqW�w��fD`���$� �O"�2|�x�'�{��|�t3�e���S2�>��,+$\�M��ࣣ�{
��lҷgᗄ�xl��]���ҏ$ ~x==u�l��~	��c'PV�����[�'��#��ee[V	Q���7�5�h�5,Wluϛ�?udF���ˏ��Z���G�dE�h�����RyX�K{�(U4��\r�<Uee���R�}vJ^��u�*��?�d���&���}�7�v�k]m��7���
�Gbh��,������0��/������-Ӥ�v��د�r�QA�ј�;-;*�7�����G3҇
I��)���W�w��fD�Ɔ ���:U����w�R���y��E ��M�ee[V	Q��W< �mP�9ǧjK�|�� �2*�,��M���HaU$kX��@�?J`�p1��^���f��5��܊�W�-�4pm�|2;$�JأͽgF"?h�5,Wl�/�O'�=��#W�U���1��^���f��5��܊�iA'R�	�)l8�u0�P"G�wk����xC�(������Q�N��	�Ȓ��1��p3I��P`�k�)V��B�1/�����ٗ���3����,�ǰ��#x$E�ee[V	Q����de�ݤ��|�D+��V��m�̖˄��O�]�0=�f�U����*@mj�)�G�O\f��,+��(Pd��'�\#�5�'���I���y�c)�h�<om����4�&����Z�׍�R��ƿ;W ��.���:�Nz�]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^�d�@���G�M��hb�Nҷ`=�}�Vݨ�W��]���uc��̄T�٥��TУ��xۛ�>�u��8�x�iH3�=���B���ꡝ���#RuZ��D�"����DZ�NU�=��1�������g�Z��3��a���!@�f")u��r��܌;���'����u��r��#�աl����aGl�97��EN�y�JB���PY~�y����o)�T*�c�Q��Ne<��t��7 �E�!6\|����?��������J*�Rs�08�b(����:����
�ݚ�Н���te�*EB�̟�1J�	�LÆ���#����-/a8!�`�(i3���8�2����o�W��g��Ȋ�>�������Ra])n#���r������{$@d�̟�1���	���#!�`�(i3�5ߧE4��9�d�L��d�@���G-*��j�J�	�LÆ���#����-/a8!�`�(i3���8�2N5�Hɫ'���+m�ol��Ә�~1S�vw�b!�`�(i3��jVѭ@!�`�(i3��i��}�12�mj�{�N<'��I!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍu���q�_/;W ��.���)�2�r;��|BL˓ }4o�X�G[��l÷{H�D�d�@���G��3v�qnQ�rVY���K*�O���t�h���rg���̟�1�w�H�-4b��he=��$M��J���]�Yl;��|B�A�ω�K��� �R�QبM��u!/��"�*�����M���R��ӟ-���4�&����Z��hs������No�ߏ�����"?��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv��ߎ ��E�5���u�L���nF���<�W�.�P��c3��4br��yO{��`�
n��>�my$�N��]流�>���ݤ�E��p�����-i�q ���$5�nc�Gy=��g����Ǵ=q@L����F��� ��f�{_8�Y��=�}�VݨuN�wAB��O���&z�вԺL�9�T�I����y���c��ᥟB�'��a�S���%�����ռt
�AԢ�a\蟟Q��ǺΕR��ӟ-�q�x�~<��w���	�e�<j��.#՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r��;�jmT�#�YN
��)e���^b�~H����8�O�5���1tSjv�!�`�(i3�YN
��)e������p�r~�h��ݚ�Н���w�w:�!�`�(i3%Q�[�J����˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 ��H�����4br��>�=,W�[�?�R��n}�����Hٚ�-����!�`�(i3	�)��&ghRV��R�4br���h�Һ�!�`�(i3��jVѭ@!�`�(i3	�)��&ghRV��RK7͍��|��W&":�ݚ�Н�$f��_Ub���r�������W��{��I�+��X��WG ��hw�U�1S���%��V�c���Ǵc�1�RG�p�P�m��������a-6�DaA�іx�~=&lL�i ����yw�kkr��;���};#P�j2E�?��˓#����j�V܎L��dE��İ���K7͍��|��W&":�xȀ��D׏�����Mp�-a�D͢q��`�L�x�$�M���)���߄�	�\M?��y���L�ΪA��YN
��)e�*8Җ�N��k�=H����8�O�5���n
V~$�j�V܎L������ⰷ���4br��$��x�-O��T���B�R���>_��\��;}{�t���=�gdN�<@Iv��nt=:�z�X
3kZ�x(�i��/R�P�HS|�O�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�k��{`.~��No�ߏ��T�4(���;��|BJ�U�� �X�G[�wE�=p���4br����3v�qh�5,Wlr�r%)cAQ17�b�����d���!i�/��mS%rƂ�o��+rp�叧���5ʦ���'�QV[1��<[��a�D��<F��� ��f�{_8�Y��=�}�Vݨh��J)7�������<�02r��dN�<@Iv��nt=:���/z*x�n;��|Bʦ?�H#F`�� �R�ćTm���j��u�Nb#¯��TG6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r�������i҆�w��kf�6�(�A?'���c�e�|E��΢�Mr��p�ԍ�S��4$:��{K·��ΥT�tE�ŀ�sb�*� �XU�*��l�lG�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�� U�9��n	-�L��&PY~�y����o)�T*�c���&����ŷ�k��d䖬n���S滑����ZLN�	���:����
�K:+>�͵�p۱e��0���J*�Rs�08�b(��MdGN���!�`�(i3�a;���a��Bf���͵�p����#�=3!�`�(i3��˓#��͚��m�Bx&����˦G�����"�fĉ>99��A0ok��fĉ>99��o|k�Lb�"������U�._�h�5,Wlr�r%)cAH�Ћ�r�H�RtV�^�G:w��-6�$�Dr��c<.~\�H��/Sg�w��'o�MdGN���!�`�(i3
x�ߜ�BɆJӱ�zW,D#kZ_�U2����}Dq�f��	��x���"n�Κ�-6�$�Da��Q����ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�Sm�6��`4�04�jf�*4��%�#o�]�ʄ�	�)�N�O�W;D�0gv�%Z?�R��n}�����H�-M�O��~��rpf�2&tRW��n
}vh�xC��f0� �-:���h��e�z����,_�k������I�3���o��(fw���'�̗������O�j�v�Ut�\�� ����%��>M����?"3�m�����h�n*��(� �C� �1�����Ǹ���)/�~�T���]�q9+t�}8BW�R7���r_��m>f��8�D�u��u���)������x�ԉ�>x(�i��/R&����1㋾����IdN�^�%��>M��_L�"����A|�stUy��{oFU�b�$��Ut�\�� ����%��>M��_L�"����A|�stUy��{o@�f�WfTUt�\�2b���J����w_���!�b[�Mv!���xB�R���>_��.�2��0tNF5��q���v�{n��뾦�c�}���Fo|k�Lbx(�i��/R�;b�-�2�׏�����M�[�S�n�H�,l����M?��y��W)�x�F[�-6�$�DK�(+�`W��,8���|b�,�ۮAH�œ%�	�)�N�	-�L��&PY~�y����o)�T*�c�p��;�{��,"�~�K���9��4�Ä/�,o� �ҋ�;��.�[ ٓ���p��e�_y.O�%T��C�~0ޭ�A|�stUy��DbY}n��!g�θ�8���d�W�J��H����8�(����X��WG ���4O/3�L�3B�\G��C.mg��n��뾦�p�-a�D͢q��`�L�N�]�B���vE���GFOg�S�<�c�!���X���z�`�|e�3B�\GJ�8;��w�h��Jc'�yK�w���"X��[��Q[R�7HN��R��bP�63Z�t�5ߧE4��Fr��jCZ�zk��X���#7�I�Jw��3�HU6�0�\��S��4$��}���`�|e�3B�\GJ�8;��w�h��Jc'�yK�w��
��Q�# 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��Wv�A����w�V�"~�ӵ(r7�8� ��$d������`7�tȈ������9P�-�,�AG�<���X饿��!�iv�aQ�Ϧ�M�ኾ���L��r�U���f��/?L���u�D��D1��n������� �k,
"i�̄�ѭ���ɿ�kF��l�l"��l䋬5Kq!�`�(i3!�`�(i3}��[b:��'(K�lc���97PC�e>2Tg�չ���1Y]H]w�
��P��*|��P�˩eNUD60L����q�?T���T��� ��?c�ĭႿ��h�q��r����$l�
�H�t���� *ί�$�E�#s�ss�7\�	�������;"��*G�e[u�;0�쒕��l\�����=@��Ù��\�����;��c���X��3i�+� a⣃_B�M�˵·�ۥ�Y�m�չ���1�]����7��j���N66j�"HsplS'yJ�p��)�}� ���x®�{9�%��t���8����Z��zH��\NیL_��f�Ä/�,o썀���P�e[u�;0��?w����3�s�'��U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�JnFݲ��s�5�>U�m�j*��{�%L_��f�����,���R�e�0����[�4�f,�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r���s�Yls��8��GM��-����!�`�(i3����]dF!�O+�|/������Lx�A�B��8�nb �z�g��U-�ew���7VaN�\�]
��s�G��38����]dF!�O+�|�����˨g��U-�e�,���6+�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��R_�����xZ;a{-�X���!1B�0�/N�\�]
��s�G��38����]dF!�O+�|�ι�l�-䤔���8@[�_zβrE��g�Hbw���1����*����OE�)�%E��'Z*)�?�R��n��h
:h����t�h��W+��W��*#�m z����Z��oE�g�������(ӈ�����$��LSm�f�e8�1ޞ��&e[u�;0�2����k���RN�-#���$�m�7Y'��k���=R��Ԗ�A$�P������5d�C#/<���q{y����i�q,?5q��7���9��e���W� �{Z+ճpo守�ubs��2[�a��o���H�RtV�^�<��	B�ɔ9Q<ϯ)P<�ܓ�Y�� л�����g�Z��3��a���!@�f")u��r��;�E����=�O�-v�*_�mS8<�n�ݚ�Н�@20߀�����P0����3��x�p��!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I�Ɨy�"c�|����"�`��P��*|C#/<���qL��M����4�	��������A$�P������5d�C#/<���q{y����i�q,?5q�+�#4��F��8M�� л��'ž1�|�'����u��r���G��^���J��sr�lE�g�������(ӈ���m�r����I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^R���Xc��Yu�����a��� vc�jj&��G�9m6�XƤ5_���"~6���aq���s{�'!�u��r��<�6�Q=2VP��Ѣ��P@JɈ.���3R��6 y2��R�\ Nh�;�P�t�5�� л��5ߧE4�흔\ Nh$�)�vx'X���5����'G�+p�9���?�(�JZ�Vk�;��|B��loXBȱg�S>X;Z�˯��R����e���Wƍ ٻ�l���M���R��ӟ-���4�&����Z��W�\7�(�ɔ9Q<ϯ���쨷	
P���ɒ�!�6UVo��`�m�;����^F�=�_�7V�o��_�Rv�䩲$����tb���~�26��\� :����JHn��z��r9�3C>��Ӛ��S�J\7CZ�zk��X��z�1P�үle�0��|#HK��A(�c���_G��Hb� h�ҩ�pi�NWHC�ۥ�Y�m/��kOT�����y������	SN��r�J��p��b���Nq#5z�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3�#}�{��~v� 1��&k@C�Ɨ0z�cULE��K3�jAԢ�a\��ĂB/�缍kv޶Gla��Mp��֙l@�B�!�`�(i3�kv޶Gl���lr�q��p��b��������/!�`�(i3t�td���5;�jmT�#ʬw�S���d��-��!��EJ��7ޅ7�=w�'�̗����S]�_�_��u��r��!�`�(i3Sm�f�e�=�⳿P��}Dq�f���.J7h��,?��&�)�
�k\�i��}Dq�f��߆�p�h��{$�������LQ�/8۶&��L�H�W�J��H����8�O�5���1tSjv�!�`�(i3�Н��Ei1.��2����|e"�B�'��a���� Ev��\��;�,
�:qEp'{w#/ B!�`�(i3Sm�f�e8�1ޞ��&e[u�;0�2����k��d����j��8�u��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��}�6�nq�Z�@���v0��L�r:�}�6�nq�4�	��������A$�P������5d�C#/<���q{y����i�q,?5q�+�#4��F��8M�� л��'ž1�|�'����u��r���G��^���J��sr�lE�g�������(ӈ���m�r����I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^R���Xc��Yu�����a��� vc�jjM�ｂ g�����j��8!��?V0D�	�I���_
�u�Y���H�hbvk~�#x�DS�AvF̓@?5�#j�o���&�2��������j���L�F.0D�	�I���_
�u�����|�G�p�P�C������H8Џ�Ӿ���yi�1tSjv����y��lD(�D �6�|�;�ƇT��J��sr�l�ԝy'��� л��5ߧE4��<�6�Q=���F��O�C#/<���q��ܐ�}ī:f����p��'G�+p�9���?�����,�ǰ����adp��e���Wƭ(n6eF�/�B|0<2��'7�u
f�.�c�n��`�7�,��n6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�H{���<�e��BFbs��2[�a��o���H�RtV�^+���G����$�\%e��}Dq�f�#� �,W���Ǉ�y!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^i��H�p¢	�B�d���%������4s����ڕ3��t�ƍd��U>�Q�c6��?��!�6ʬw�S����}Dq�f��5ߧE4��"T^r��~����k�_�mS8<�nZ�~�|}�"����Ż�&ǥ��bP�63Z�t�5ߧE4��Fr��j��k���;V�
pFV�$=+R�˩��*��� ��U�_:�E��t?����a렾����޴8"��J�a$�Y �t/�(�P�KZ	��\#�Z¥���5.'MtZ�R����DZ��}�1U��VP\@Ww6CE!H^��Ƨ�0/��U��|:��'!�P�P2����+�wձ}���8y�����e�Q�� �)ԴG<�鶰.����܍ \O~��z����
����7,������Z�ך�>1Y�>c��?�B�t�xr�t��b����J�"I �����w���'�(�]�[�H���,&ǚ���φ��<�6�@a� ��fFMqlg��z?F�#��S�J\7O.�x�����(���2$�m�����G�'ž1�|�'����u��r��RD�~���M��V!�D��nF���<�W�.�P�	��
�Q�}g��A�L��d��JXl'�T��~��Uг�|<m�����G܌;���'����u��r�����Fz���2�b=���i�Wg�l���鯻��U��O�D mWNs_ѧ�p�O�D mWN���J�a��IX0F�Mb�Xϋ?@�n���/l�̬���	p|�O�E/�9��"J j�E��'Z*)�?�R��nj��P_Q����t�h��W+��W����uR���_�#g� |cz�����]X����7�4��~n�2o� �2�L2��R�͢��n-΂��m9Ϲ��*��x��� ���JH����8��#I�ND�s���H�V��-���^S��$�Gy��e���W������)<��U��)���Y;e�iK!���d."�9ŭ,iI9�o«IX0F�M��ŊPTWo9���b��|2;�E����A(�c���_G��Hb� h�ҩ�� ͷ�	���6�
V����b+}y[<�6�Q=�B -�6���'�QDndN�<@Iv��nt=:��:5A��p,�u�S��d��JXl'�T��~��Uг�|<!�`�(i3���9���LQ�/81tSjv����y��lD�TaDe��"�/֖�Yk{:fh�3�:5A��p�� л���������Z¥���5.'MtZ�R�!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I����~�Lk݁ 1���tw�i�Ք�w��y����J�a��?�d���&�J2���n�7�ct�����?
Z+6/Ahr����B�z���b�~8GJ8��"'���xO��H{��4-�9���{��Psmi'l:}��Q\�>�7���o��_�Rv�䩲$��V���,�wO0 zK<U|r���3fX�?���'��>��ԑ�%;�E����A(�c���_G��Hb� h�ҩ�h�x��JyW$q(W���ƍ2���l��^{T~H���^a�nu4Bޗ��jw�	���ݚ�Н���fCI��8��GMZ���Ӗ���mFA�$�!�`�(i3����,Ů�뒒���97��EN�fԯA&b닓.�`�3u���# �%��,�V�B�
X��Z����b�Ի�!�`�(i3�(��p�m���
y������Ľ���ANʂ'�8���y}	�'C�R7 �E�!6\
��7t��i��E�y�H�RtV�^߇�\���*���H��w�u�M�Һ����1)uם�!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I�Ɨy�"c���? 6����,�ǰx͝�I��D�X�����t<�NA��qޠ	S�uimK�ֶ����6�o8:4�I���c�90��6:����+�^n=\f�5>�I!�[�������QQ��B�"}��r$ɓǃl[�Ƶ�1tSjv���R�?�Γ�]#�y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�S�#p���zՠ�����˦G�K7͍��|��W&":C#/<���q����g�Z��3��a���!@�f")u��r��R���Xc��Yu�������&G���y��lD���j��z$��
�5L��m}I������jH�2�s��� H���Y�����&G!�`�(i3�r���Ipˏ-).^QQBպW � ����i9v�I��`j!�`�(i3��&.��8�F�S�1 ��po守�uQw�$��Z��/�dW���3����V$=�b�oj�+p�K�J�iN�Sˇ^�6�H����8��� I���\�b��v݋N�����i�!w���p��;�{��!�`�(i3�<��	B��D厺��+�̟�14�����{��O?��ʔ��,Vr<�6�Q=��jVѭ@!�`�(i3S�#p���zՠ�����˦G�K7͍��|��W&":�ݚ�Н�烉s)�v�bP�63Z�t��Qѳ$G��A0ok��烉s)�v�T����� Ԕ׹�Ӫ��*$���A�<M��[��k�}�t��/�dW�<龈��ơlП���V03Y��9�`�I��W����Ľ��M�ȅõ����(�x�HM���#g�s�
�`�I��W�^��D����jVѭ@���Fz�!�`�(i3!�`�(i3S`�@�4:��]�����n�h��N�M��~��f�!���zՠ�~��q6g�yF}���V6l;�<��'�̗����#!d�+I0���ԏ�.fOe	�N:w�h?Y�)�}���"���d����yi�l,V�,k� sȸ�"rR!�`�(i3�����z�>9G`�(���'�5�,�xs�*"1���)�=�w�������:�5}`'l:}��Qb!��u����$A�O1�Et�]�!����M[��Ǣs��j�ŉ��m�n�~�!�G���-7s�9���o>��l%i�-�F*D@��j�i�p��+��~���O!��Q]� _ό���.��|�����E ����7dh�?зq8�Ј'���Xw�,bxqX�b!��u�<�`A��_i3i 
�c��]�!����M[��Ǣs��j�ŉ�|�w��DK����$���7s�9���o>��l%i�-�F*D@��j�i�p��+�/s�1��p��Q]� _�rs�i���`�M�	=̞��>��3
�v�v-}�	mp,��_А#�<om��F`���G���`y���C#/<���q�5����`KiW��
�!C� �u؅��FJ��gm?2�I��6�]���~`��ʿ��^�����èV�H�?���E�m ��?Z��G.�w�v�d����x�l��1:�N�*�x�� л���D��������m#p�W��	]�	M$E�Z�ݚ�Н����iYM�5q{! l��2
L./;�Ly�Af�?ǉ�=񔿄�aB6Э~���V��2
L.�X;p`��3
�v�v-}�	mp,��_А#�<om���'$W$�X�<�6�Q=�L�K��%<7�`+Al��R��������,NL ���<�6�Q=�o�f�Ԝe���b�!�`�(i3�(�;\��B�}�ݚ�Н��D���R]���gRI/!�`�(i3X&|a�#g()��ikp���H������7Pr��ġ��,�&�C�/�s�f�I��b��v�#$�q�
k-���w�E�V{�!�`�(i3�V�����/>�"�Ax!�`�(i3��3�N;C�]�'!�`�(i3�7Z.m�w��'�k�f!�`�(i3�u~xgA���������6%�a�k���n�}�� �с�'(�U�c�&8�,��
�Q!}-[BvGޣkQ�A���ۖ$����nQ�rV,?�����ݚ�Н��43S�d��ރ;�{��C�{����K�7��C4%̈́��� л�6�R�W� W��|E�q��w\F�M$E�Z�ݚ�Н�H���!�>�*�!�`�(i3���K�7��8C+a�Rj�~���0ȓM�Me��^��>�z'�:�N�*�x�� л� ��$�,���X;p`����$AA�:JϮ����j���ӱ}�tM�@;w�$C,0�?���<�6�Q=4?s����k-����b=�<�6�Q=�0V32;5�-�����4)cq�vG+|�<�� л����ٜ�]�X;p`���C�,�4���y��lD�Vf�`H�j��-@��ey�E���x�ր�ݚ�Н��y�3���k�K��hczZ����4b�zvѓ�!�`�(i3�7?�S�!!�`�(i3�$�~c/~�O��������y��lD�Vf�`H�jT��b9���ey�E�����$���f�?ǉ�=A#�
�v!�`�(i3��%ў׫=�F�K�@�!�`�(i3V��uL$��!�`�(i3�$�~c/v��&EA)�� л�֕ߝԀ�#kcBTX�#�
�ge[I��4�	����������P�=��:F�|���m�:�-22�v ,��rQd->�d�!�`�(i3f�������9�|Nb��'1-�,bxqX��ƿ�d���5�[՚1D��c�e��o����B��7dh�?��,:&���z2%警�d��]�Q��f�_��BvGޣkQ�A���ۖ$����nQ�rV�}!�@�?0d׻zc��7U�	Y���۠ql��*O��_^=�/Jt\�J���70�'���O�V2y/�ߓ��y��]��K��Xw�e60�' ��[w�{0
����)��#L����?;����IX0F�MV�ҁGG`5:��0}}��*ꅺS�J\7�p���"Z�v��!<�6�Q=�r$ɓǃl[�Ƶ�1tSjv��� л��	�%1A��b+}y[��\ Nhk+Q�h'�Ȝx�5W ��̫(� h�ҩγpo守�u��"����G��Hb� h�ҩή� л��	�%1A�qo<�khku��J�>�V����f�z��SR:g()��ikp���H������7Pr��ġ��,�i�/Q�ಧ�y��lD&[�x�R�"��}Dq�f���&.��8�}Q�sd��]� )�+��p���"��NwK�"&'��Y_�C#/<���qH^��Ƨ�0	�Ʊ�R���uoJ`AP�n�M�t䖬n���S滑����ZLN�	���<~=��<��?6Ґ�6�d45sf��ݚ�Н�<�6�Q=��b+}y[R��X鷴QW�w��fD!J��/٣׆p�9��+:��0	��