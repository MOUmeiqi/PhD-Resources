��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:��ښ�1oM�U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]���<�j�C��`��L&`^����8��U�Z봣��D��L���_�L�3��0I}.�ANMs����Ѡ�/�Ҷb��N�w	*D���y&�f��+K��[y��ڂj�x�z:I(wKq���/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�0k�5k��J�|(���u����l�|���j�I�?g�f��#��� �bRw�����IL�+�{Dr[��=�^S���Z���y�ۘ�G�|0$��&�^C����Jw�)��Pip<ɯ�nefR#O,.�c�u��QF}����;�A3�'���/�k��±'�R��;L$]��]{�[N�4�=,����Ϙ�Ԕ'�Ӝ[Y NoC��c�S+d?S�7�$�>Y9w0�R<�CW���V��r:O!�`�(i3�g���}���������8*��#�N��O���:�9`�p�0��&�����¶	�Ev!�`�(i3!�`�(i3��1�<����>l�ݯ���9��)����6q����"� _�i��i���5���6*�t��L�kjt���?�����Jm�W���K���v�7��٤cF�Vq	�!�`�(i3!�`�(i37p�J��PW���3���D���o�i2��0�ּ���)��G�������ϲ���>h�c}����>I	���(��B�:����@���4W�-c8��"�a�O>*�ׇӭ��!�`�(i3!�`�(i30R��=	�@����W��nl@O4茸z���q����R��C���CS�� ��!�`�(i3!�`�(i3�0�9&،EB����n��|1�b�YL��&\VI`,xJ�����gc �{�=2���p�)U!�`�(i3!�`�(i3X�o|3����x�u��"��휺�&\VI`, �DO'�L5я�����0��zO�)v��$�Pr`7ï&��.�-�&��4�%�@V����S�����Ŀ"���J���>�$!�`�(i3!�`�(i3H������gf���5��x��X�mϒ����y��f������E\/P*i��!�`�(i3!�`�(i3!�`�(i3 ?[n�:#G� �b�H~V�I>1͊���3-���I T�+����̵��8<=!�`�(i3!�`�(i3!�`�(i3C �@nk�@���;)�����<j���ֵ�Ů�y��ͮ5��}��6�8�-Zy?X�`:;��
c��@*1�L� ;N>�G�$U��ިB�Y�5J��5:5J��(�ߜ1�ׇӭ��!�`�(i3!�`�(i3!�`�(i32g���`����&\VI`,J����^��f�������W�� �!�`�(i3!�`�(i3&��潹��a}	/ȸG�$U���pJ`��8������O�w�V
�1!�`�(i3!�`�(i3!�`�(i3�I��(,�a]�l4���?�AO�]X��ƞ2�� u8�"�6���G��ꚕ�(q!�`�(i3!�`�(i3�EH�2�L@���_r�Gl��c��#
Q�����zwK35���h�w�)ꣴ?���X�!JFh�`������eC����	F�o�=��KQb�KK�y؄@�!�`�(i3!�`�(i3`RXK:�w� 1ܮ��gf����;��@B�a����K/tE@��j�g��o��,�r8ЧڜX��hvծަ� �0���o���Ѯd.�6��S�6�0RD��}��b.զjUǡ�9�ă@���3)ͰnL
sȸ�"rR!�`�(i3!�`�(i3�z�:>�=��9�V��r�-b0��[��u�j��-xIYBN~x~,[ӝ60��,o�!�`�(i3!�`�(i3!�`�(i3Eu^Q��X�[�"�k�fQ�����z�xO��̋z�:pF��w�=���6�t�qŻ
p�!�`�(i3!�`�(i3!�`�(i3k��U_���nཱ�&������!�؟�r�Y�}94�h	U����f�7U�i�#!����P�>+�va��2	p���>/:ܝ	�@�ׇӭ��!�`�(i3!�`�(i3�>L���L�ɚ5���x�[�%���%���=���pw�ۢ2��vR�J���}���	��!�`�(i3!�`�(i3����N����������(��K.���ccnh?��7>�����D/͘B���&,��*eM�����3�j��~[�h��\�ڰ���gLE�z�K�y؄@�!�`�(i3!�`�(i3�>?v��B{?a� ~>J*�ya(�$>&�.Q%�i
u����-1<@GŚ�ׇӭ��!�`�(i3!�`�(i3eI �#��I_h�R$:7��}�؝�T�D24N<I8����\.Wֵ*&E�^8��xt��:_/�~8����A�߲wLB�w���#✲�@�킍�"�?���Fz�!�`�(i3!�`�(i3�s�cn0�u�A�qL��D24N<I8����\.W~C*B Ɣ��(J�fŊJgSᚄ�j
��a��ǂK�O)��+`�{�gt�R2���4eM����;�0Z�8��1	/��R2ռ~�S�N�\�:����{����~��➛����Xw�e60���Ϧ�lـ��Z�>�=��$��6��{ֱ@���O���:R� -�*3fх�-�@���q�qp�HTEn����1��7��w׸[�	�+%�����;�e >�#�mi��,�kL���Pv�����'Q�@RͤUʐ�{?a� ~>�8�<��{�#:B�6��1��h浏��������S����3|��@$�g�9f�oF�7�8��i�c�������7>�����D/͘B��)gI�qd��+L{��+x⣗�C�|�6G�"	�WJ�Slm���`�7^�	���*�C ��s�Ε?�������4��A�Ww�=�d2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hͥ<#���vSB��n
HDW�Gj��o�/��];Lth� �K��G������\ͬ�W����]��Q��S
�yl}Vİ�M�W9�f^�Ԫ^��rL���	��D9�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc	���[�;�4A�B�'���W����+n2Xh?J�k;��7
��t^�L3��헙��l���Cf�O�P,&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q��f�SR�v�����������\͜��ͱ�5�����\�� �K��G������\����h:�Ê�����\�$90�H1�����\�P��y40�^�����\�T��v�`2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������w'��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:��ښ�1oM�U���T�����\�4�sƐ�hd	�ѯ������(�1��_�H�X~�P79Ř��W(�̽^�T����U�E�0��5�Y�w���ؤƂ��l���]����?�AO�] �\Yy���y7>�?�}����eպ�#6M0��I��7�O�.$��Y+1���u�#��ntEB����D��;��M6<���gl+�����p.;��|BG���pi�A9��g�L/��@3`K�%u4�+lnwG",����
� �AH�P����w'm'���h$��ޝ�~J�'v���"�F@�4%�}����b�+gobQ�el���V4zm�!=�y����h�}��/A�#��0�.�	�Z�����}�P�y����E��Gw��f c$����X�KM�^~$0��{�6�x*�R��=e	6'��}xYϷ���x<]�`Ý�M���A�t�>�c����P��RL�a)r��fI�������i�9�0NE��y ���fνw�>��S�@~�w��!+3��n�-��U��N{K�s���ʷ����# �u��.t��3�`|�}X�m����D��`7o�����Ѝ���z޷������RL�a)r��fI����D�-��9�0NE��l� ���3�w�>��S�@~�w��!+3��n�-��U��N{K�s���ʷ����# �u��.t��3�`|�}X�m����D��`7o�����Ѝ���z޷������RL�a)r��fI�����,�%��/w�����.B
'����u���;� ��!��_+�8�X��m���l��"��QpR6P�?��ԭg �s�~�R�3ԭ)&l�d�c��t�jPP�
� �AH�T�t��3�2w���$�c����d�r~eIµ�Apv)!����e������~C\{��RL�a)�O��u���I�~�CVBK�qX@oXeL��!�zg�Z�$����O�V�[1�7��s�M�pD<�x�?d���6С���^3��/���m�!=�y����h�}�)��� �A�s�j���2tt����Sd,�ϱ�ϖe��!����i�kJ��x�l�e���#
��� �� �6���{9�6�k�8���҆�|n����vJ�^1B�f�l�Z:K�`�&�ѕ���`����/�~8��Խ�Z�$e�246��pa�\�(Xc���0ٺq�s�ݝ����vȯq��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�=W�֯�ZW���xF���慼|~09h�i�;���6�ӫ� n[)Z�Μ._^��/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_/����E�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcd����ɚ
	���qk�ZV"���:��#tC������s�F6��UQk�!���.��e)�Op$�����8�#����S��������Ǜ岦�%I^��������D	��U�e�n�^��]��g3������ɤ|pW�Cy�w=�4e=��-��ؽ7$�	�s}��[�wH�HͶ���ܜ?n昼�2#:��b9���P9b��	�Y���1��� �U��֜��3JHn��z�C�$��؍��R��j�.(Wx*�_F�k-�!�`�(i3��|g�Y�'���Xw�������펎��{5Yl���#��]���>����Cί0C��؆Q>�[G�-X�@�^��1�(R\֎u���sRt�7G#+��\w��0](@X~�H:�W��7=c��Et��q���U�[��N���v�Z�]2�y�Z鎬�����	�7 �#�\1^O��0ˋ��I��w��,>����C��(R\֎u��ԟ'�D�7G#+�Ǘ0z�cULy`�_I�v��4���OTWRdr�Jbk-����'�\�n�wa��>���g��U-�e�,���6+�=�B4˖ב����E��@IE�U��*�QN��� ]���f�fx��V$�w�I�?g�f���\X�<����8��UWJ��)��q鋴�*Х�]��:2�R�W�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcq�P ڨ�| c�]h�۟�r�@m��+�<4��ˌ�ň��h��j�V��vUQ�i��7��!�Ԣ��:����@����gG=%� g�Vv�5)��Z^7s�9���o>��l%i�-5�e`��9�\1^O�cɴɫݜ�Z鎬������_�,�[/�cWM��@EZ������Q]� _ό���.��dŚ1N套�qD0�L�I��W+`�x�o� E�����(J�f�6��Rq���8���/��n(���˧�0z�cULy`�_I�v�1��� �U��֜��3,0=]^	�&|#9���b!��u�:�HCaIMl�=��套�qD0�f��p&dQ$n�ti; �L�q�t�MyފVZ鎬�������(���"c'��ɿ���1T�XQ/)�EY���������S8��>,�����$�Qu��
Uc�v7�i3<�f�D.`�Z���N}�m��{A8�#�;:�H>+�w��0z�cULy`�_I�v�1��� �U��֜��3��"X��[��Q[R�7N}�m��{;ڋK�m���n`5�fK��0z�cUL����!�F�8���/��8&���IS�T"�IÉ<i�LE� R�g��U-�e���\m�>H�)����Yk����B�=����g;8�ݚ�Н�޼���"f���Z���{�u1H3�K7͍��|��W&":�ݚ�Н�v�ܽ�oԃ��Z���{�u1H3�O���嫑�!�`�(i3Q�#��݌Q��������$t���$`E��Ե��6���f��t����D�muշ!Rq4���u�@9 Jܵݓ�W���2��lKA#ݠ�m��/N+0�-zNvj)����r^ʁ���Mյo��6Z�L?��:�پg�+���C&��G�&ց�*�+��d��h�6�q��� �pkf��8���&�(*�O�q����╺2N�3u�&��|������}Dq�f��x����իU��j�/T�<�_�y&��S�ݚ�Н��gv)z���Z���{�u1H3�;�У�M�!�`�(i3�J*�=[ǿ�������$t����]䍤J���6��J�|�-&/k�D�mu�#��bE���u�@9 Jܵݓ�W���</#^9wlݠ�m��/���%��ōj)����r^ʁ���Mյ�����1,�L?��:m1<0� 4M��C&��G�&ց�*涼0�H[��h�6�q��S��"��k�8���&�(*�O�q<}��kUEx��2N�3u�vs��?����}Dq�f����'��@�my$�N�j�/T�<�_k'Ͼ��;b�-�2��Q�������|#HK��ze�9Up�rP��OA�/C��?����\��_Q��ڋj֓�D�l�Q^�MY:�H 䴢��H�RtV�^?#1���2��i��>Y+ѕkOo�~�K�$����@�І�y�!�`�(i3!�`�(i3!�`�(i3���b�3!^�3�@ym��[jpe���#׷�`�:\�Q^�MY:�~��;�,�/��@�������̠sxd�li?��t�uJ|���8�� ���&l[�]h9��`y����;b�-�2�'{w#/ Bl�i�<�9BpS��x�f@��S��,�����`�|�XCtK[j*�4����Ě����E�i�m}640�RS���$
�)R�@�6�֐�2$%-��%sEW�o���開������
�9ze�u��S8�RU��E�{y����x��F�U| c�]hn���Wa���'(��S1�ӿ�Q���'(��n�FJ�>��\1^O��[�~�����\1^O����^����0��G"��������0��G�ΠE�n�m�j��A�7�]X]����,�\� ��%�D�v�l�Ū�TD����>�֔،��t�h��W+��W��7�]X]�}�4��d��D24N<I8����\.W^�V]��}���_j�Nh�EC��Q^�MY:�́# (�套�qD0Sh�Qc��/z*x�n;��|B[�x��ޗg�%���۞~��3R7�j�8`�z.1�1�N���PϾU4T k���%f/MR�V��Q+��
���:���
W�&��9Ԍ�����!�`�(i3$H#Ö�U���KX}�!���ra�[�k(���"H�@�өN}�m��{�K|��C9*�¢ڎ�����:i.ߋg���~�26��\��%�����d��9�ՓN5Χ��F6l8���x�;���EWr�i���b�Ȇ�� H�qo�:�ȧ2N��n��9:!T+} �f70���"�,�>E��ʆ�In��t��+x�r�s�*�IŰ��� �!�`�(i37�ܥ��2�{�*L����Q^�MY:Z��s��u*w�A�2N��n��t�J�Yy� ׿`Hڛ?A����cforS�b�8Z���oگ��r���%��Q^�MY:8<�a���D�P�E6����{�d=��¾ȼ�Zj���
Owgn��ݫ�񬿱U�׉YH�$Yu��r���5j����b+}y[�wbk�$T��8$2OU�1Q�\��^����;�jmT�#�	�"O���V=}�G�����&G���y��lD��2SB�tᚕPH�ZØy��j��k
�X�nZ����}b��:5A��p� ͷ�	�"Rc@TahbIQ)vl.-����a�~9��tf��!Z鎬�������$�y��j��k펎��{5,�Lǫ�>a!~�)�=5U�i�J�8�7���}Dq�f��q�	��c�.�h�x�~�%!���wbk�$����$���]�!������G��+�t2�|�;�Ojz�!��_�*9 �$R��j�^��ݔY�{'%suE9�+����Q�Y�<���%�� ��0d7�y��j��k
�X�nZ�>��Hh�Nyλ������ݚ�Н����L2yP��C��?^<����3>a!~�)�=5U�i�J�8�7��S�Ĕ�Z�����'?�5�o��K�W����E1��a@����}��c��v�q	����7c�	^�+��J@�h�����XX�<�6�Q=�a�W'������PV��y��j��k
�X�nZ�>��Hh�Nyλ������ݚ�Н��(R\֎u����>^17��$R��j�^��ݔY�{'%suE9�+����Q�Y�<���%���!X�I�Y�wbk�$����$���]�!������G��+�t2��\1^O���)�`�>a!~�)�=5U�i�J�8�7���}Dq�f��q�	��cE}k��9�O��F�`,9�H�W�I,�D�y:#9�]�B�_��wBW�MM
��,=*A&-�Ri���y��lD���|�D+y-ʲ�}!�`�(i3�;;����)��U'���>
A��%���ؽ7$�	�s}��[��-����!�`�(i3T�8o��7�Ft�[���!�`_q�!�`�(i3EOJ�uxm�PQ%cp��g��51�X�c�rs�i�}�O��LTSG��ʎ���d,�0˝Sz��E�4.@��n��I
�:qEp<�@b`��%R�W"���z�X@*[�]�ʭB�?�`u��r��!�`�(i3~�`cC�4��L?��.��� ׿`HڛuE9�+��!�`�(i3��܁�c��ލ]	���{��mj���rs�i������%!�`�(i3w�����A��ߎ�x��yW���5�kX����3>'���Xw�j�7����NWJ�2{���G��#!�`�(i3\OW�:��d�}��v�%� (��Q�ce�c�Ԛ�-����!�`�(i3T�8o��7�Co7�wk����7a�YCy��}Dq�f�<�6�Q=�G�)�<`�4];ˍH��6�,��)20�	�:]If���ՆnZ�va�?g_����24������ȕ� M4x�Q?M8�f2!�`�(i3ݜ�
N#�'���-b��d9=���u��r��!�`�(i3q�\E��0N�]|-j��k��?���b+}y[!�`�(i3�	��x��ݚ�Н�!�`�(i3套�qD0�d�i��?�%�_SK���|e"!�`�(i3���F��O��ݚ�Н�fĉ>99��R�Q���~��p����
�:qEp'{w#/ B!�`�(i3�����*[wL>r~�/1��0$�������v�W~��,��=c�CuV��A�
�����=@'ѥ�fĉ>99��A0ok��fĉ>99��R�V�"�0ɕ��aR����%>�rGO�D mWN�	��x��ݚ�Н���Aj�%����NM������F��O��7�癆cgjF�ཕu�dZ#'���;�#}��\"]���sN�W���T��~���y�:�����jVѭ@$�[6{�!��N��I��t����75�\Gg�e���%>%��45���\}9�z~S������:EM����Lg��gq?�������H9��p#�7ڊ&r����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ſl �