��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�>���U�_�4�0S�����x�P��'�<7\F���r����&$9g8�M>PFWD#�z":���ӳ��_}��0w�\1����K~�j�k��� �Pq���Ɽ�Yk"1/s�\"�����p"�+ڍ�P��Ѡ�/�Ҷb��N�w	*D���y&�f��+K��[y��ڂj�x�z:I(wKq���/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\���z��<�Y��{^(�Ś��
��H,7���ZXWL�sZ�	!w���� �bRw�����IL�+�{Dr[��=�K)�*�-�>�����Ádo�dN<djY���o���F���e����n�QX�v����<.���+��T����oGo�Z�������/�)��ɖ�c�������]P*mQg�@zh�S҆�|n����Շ_ Q �Q�V䙔<�[C�
kf�+������u{Bo�#�����7��J���u��w)�S��X3����~篟|���}r�w�6��ޓTS8�:r&@P`��dpfVpb��#`^���w`q�eE�3u��g�~p!ۓZ�)����;�*z��
=z�.(��lY��_�	�� ����J��̅��1��pp���b:@������qθ�OU����EWeIq		�]H���_�	�� s�nTNAi�ΊWw
�BAW�~Di1�(q;����d��翑��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"��-h|,���(����>S��ә�����/�4�}n'���a*�x���� ����ޙB!7����ˉ�1�:�Ω�>���U�_�4�0S�����x#�x���c=Ct�z&��ÃlO ܅dh�' L� U��֜��3Y%T��BP��&��J�1�KB|1<\w¹��<d���<
DNͺi3<�f�D���X���`��wl��h�ٙ���O��Y\�J�:>���'hZ���溂�U~܎VV��EfVNN�0|]<w:�=]A��O�T=�4e=��-�ĕ|G������E���b�jT�.����$�k��WU<o^.K�}�#�J��>o��9�0u
c�Б����!�`�(i37�ܥ��2��
[���p�� +@���a
��|���\G�Y�)��Y�%�<'L�<��z��}�0z�cUL�n����4���á�~O�"j���b7|#9���[�t��#����Ea��Z鎬�������(���P����ˮ��lC��U�T�\ ��+�_0c �X�FJ�+���-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0(����!
%Z鎬�������(���`$�P.eE���lC��U�T�\ ��+�_0c �w�)��O�ҋX����>��l%i�-�M�g������{l�f|�ό���.ӳ�
�	?�<7Ê7�E�4'���XwI<��f�@O�x�7���q�©�����<�������~s���^��w|j����NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��Qө}�8o�C���7I��������q6 tɀ�Ȑr&���UYv=��8`̏��$���"���	��ע¡{T{b62�tstF�!��cܜ���,�ǰ'�J:��XD�w�п?G���7�V��i��fj�_V�VG�88�;矷m�w���i���Z��Ms�����x!)�M���r��0���u��n	l��Q;�im��ȍry��	�6�5�p���PF��W�!�`�(i3!�`�(i3-��<�ξ�\zǣ©���s�٩���I���Т��^�\!�`�(i3-��qW8+���ǣ©���s�٩���I����:�Y���!�`�(i3-��qW8+���ǣ©���s�٩���I������.V��:�!�`�(i3-��qW8+���ǣ©���s�٩���I��������|�!�`�(i3-��qW8+���ǣ©����@�hGq6��nX��U�	vn�����7Z��-�����m l�o�&�C�/�ީ�%��w�*�fBg�!�`�(i3!�`�(i3-��<�ξ�\zǣ©��
.�Ūz�/>�"�Ax!�`�(i3!�`�(i3-��S0�:�l����g�SH9��n�7�Y����Xc����L�{!�`�(i3!�`�(i3imp�7Ic;-;*�7��3z%�u�܆�=�<���XΚ��!�`�(i3!�`�(i3!�`�(i3�sg]�_�}F�r�f�t��5Z���@x��D���j�C�6̓126��G}!�`�(i3!�`�(i3ދ�������y@(8�4�!�`�(i3=���yp�.���.����!�`�(i3!�`�(i3��\��,&߰��U��f�?ǉ�=��Wʁ���p�B�E�!�`�(i3!�`�(i3�X;p`�5�8Cl8R!�`�(i3�.��Ԕ^�|n�M�!�`�(i3!�`�(i3J�]�RU�`���!�`�(i3!��I\+��M�a5��|���瀆!�`�(i3��L	�����T-��/��@������1�so��d�a���A��`�c1+��D��{<
Q ���=�Ҹ�%�� �!�`�(i3�N�v�1�c����L�{!�`�(i3!�`�(i3�$wq�����0��E|�,���6%�a����>[H����&?�!�`�(i3!�`�(i3�&8�,�I���Ut�es��O!�`�(i3�1�)�c��!�`�(i3!�`�(i3!�`�(i3�u~xgA���������6%�a����>[HNl����!�`�(i3!�`�(i3�&8�,��w�Iſ�Κes��O!�`�(i3]|If">��]~'�H!�`�(i3!�`�(i30>!j��
!�`�(i3&�2�������ȍry��	�s�٩��$�f
%}�YmC,iguq�ށ �~�g#n]E�}:����p���hy�t�]�|����*[UxG!�`�(i3�v1a{J��`����p^���XZt%��m&<�,0 ����
�n��E3���?�K?q�\E��0��A��)}�\cZ��2�!�`�(i3�%]�N����%ў׫hDG���+�/���i� �����,�ǰ'�J:��XDd?�3!�Oϟd���,��ޤ[QG�