��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�"� r����x[&gݹ��]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUPc�k�u�}�R�6�_(!��?��Xm��+���������q6N<��;��� B]�pE���	x]̃Dj#^Da����M�׍�ё�6ٕL\S��A�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω�"� r����x[&gݹ��]P*mQg�@zh�S҆�|n��?�'VX&]{���|?��?G!~Ve��v.W����(R�/3�*x>����!��?�7i9a�h���E�߀����.AC7��E]Ta��b��)�c�D�g$\�]�����u�[Ʋ���5��4]HM�Ǽ�˺�ʘ�plQ5~��*l7c,�z��T.��R��KiT��X��� -���G�zV��#�,���oJ]p�����H}C�ns)��E�$lY�G
W��V"��C���<r�<T5v�ۂ������h���h�}��b�Z���V�����`���J�8o@���q�&/�K��]X��*;o@�f��v������f�aoEX��1�T���{Q$V]���RF'�_��}7�m�!=�y����h�} ?U�B��(Zk ��U�E=�K�^U�#�57��D�[���� Ԋ�F&���͋�V��Ġ�#� ��>Y\�\$�D�|\�}��/x���f0� ��!��TN0N��\�4�sc�[�.���Zk ��U��6W��q4���D�[���� Ԋ�F&��7`s� '��:S����ք�'��-v��qK=w��#���D���i����	x]�m�Je{q�#?���/�ōy�<��=W��s�!5�&}Xa���qd��.�Yt/&W��^�,��/�Mu��w)�S��X3�����0~J���r%7d7Ө%ԋ0��>��[��F��'�`���GS��(�����s��X����?J��0�����(��'��&(cį� �������RL�a)8��Q̮�F�����p�5�p��z��QK��;H���䬙]�5�IEpԞM5PI������n��D8TLE�n�5?��蒰&^���:��a\�������n�����qz_��[�|B�����s�3�D{ud�����
>Ҙ�m�<�|M����<{���k�8���҆�|n����5��K�O����FT۾D�{-��g� ��uz|�Wm��z�h���J;_Q���Qt���~
� �AH�*��.��u� �(��B�Y�S����w�/e��i�P�GyϪ+2�Ī�>�n��`��4�� r)��}�-�0�l���jgFk�Q�l�K�c	,J���ӵl{��1���n��pEh�r�q�~�2~���RL�a)8��Q̮��,�%���=w�^B��+&�sN~O�;H���䬌��4K��l�yn�=�fZ�P���sm��\�4�si�W���
�ԟ�d ��_FJ��rˍ�Do@���q�&��|�)n��;�S�˹T-~�	�Y
� �AH�*��.�:�o�E����o!f��L��	�{�3�i�P�Gy�$�������G}��$�n'�Zvu��w)�S��X3���X�7�j�����c|LU>|G��m���>�)#i�zuZX�0a��/'83A
���RL�a)ѻtUWR����H7��7�ޑ����<��&g�7C��H��C=�)3�C����")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:I�k��S�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEAvI�AJ$1�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Q�ئS��.V&��B֥�(����5�a���V��#�x���c=Ct�z&��ÃlO ܅d��
�b�lr�r%)cA�����Y%T��BP��&��J�'����IEߺW�L�sQd�h�=3�!�`�(i3�i3<�f�D���X���`��������I7��-5�B�wj$g!�`�(i3�a�\����9�	��%
a���+P��_,��ޯ#Q �4�M�����jݭ�F���L�D��6S��X�u��
)\Y��!�`�(i3�E����F���8�TP��Vchw�D��y.y�Q\�@vs""��Fq/�bi��±�sR�{F3�_� ������,��\G�Y?�� ��}r�x�e�X�����5	���]���c�A�L'��!�a��5�%]���a(􆿳����^��$���]׽������E��@IE�U����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7��=m緒��J���W�7G#+�Ǘ0z�cULd�g>57<�C�u)�6�3A�)OqЈ�&��g3�g��U-�e�,���6+�_������"B��$I��w��,c�A�L'Qī�*pY��㶢�&-���x�'@�(��P�G�p�P�į�d��8���/������T!�G���-N�By3��<�]�!����M[��Ǣ ��$�,�������5	���]���>����C�*��^�"~H7.�;AF@IE�U��>��l%i�-]a%ڔ��E����F7G#+��\w��0]C$mQ��"�,�>E����-��%Mό���.��_F�k-�!�`�(i3c��Et��q���U�ЂDa��(o��0��7��|g�Y�'���Xw�E�i�m}6	��	Mk�rv�ј�"��Z鎬����y��|�!�p�tN2s���(����5�a���V��Eaf�#C�q�P ڨ��S���Qߵs<��7�m��+���������q6IF{b	��5����`K�i�4(��T��
4�r�%Ah�%4
>��f���T,!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�;C@����W�L�sQ��|`��'��>�4N��[���i����I��'�p�
9��x`�|��K�z��u*K6HY_���P[!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3V����(��w�K�h��q"�ـ�`���|
�P4ǲ �n�/?Sk�������[b�I�P"G�wk�١��	;q��^̽1��R��ӟ-�D�s�A6�&-���x���h;C	�T�\ ��$*��<�1AԢ�a\��ި�����|`��'��>�4N6d�dG�7:�R���Z�F�\Ȳ�r�r%)cA�%�\B�����x.�KnqQ�����IMdK�Ch��|[p2e�F;p�	+��Q��:~�G,�A@����0y�	�C�u)�6�3A�)OqЈ�&��g3�g��U-�e,%�0g��Չ3����F�x��&���ő��̼ғ�vq�\[$Q��
�̞��>���I�Ūe�TU]O�d��g��U-�ez�r�6�>��왩�>G�g�����K�M�{�0z�cULd�g>57<�C�u)�6�3A�)Oq�fhz���I�Ūeߋ٣�o{�i7�v�ԯ��Q[R�7�����bp��Tٷ��(�UtW�*X\[$Q��
�̞��>���ԜF�����`���W�L�sQ������f���[��R|#9���b!��u�̲�2�!�y��Fp����f���,(���B��ɓ�~Ҡ	��[�)�D#���ߔk�V\�5��|�~�R�wX��}�
�?����D)�ܷJ5�7��4'���Xw�j�7����w�K����+��dЧ^{�j$��XCp=8�b(��;3��o�r��`y����@����gG�G/�����<�+rAԢ�a\��F�dH�E�%<NR8�b(���sjߢiVr�r%)cA���YVO��R�wX�ո@����gG���>��;�-mO�ғ�vq�F&|S���T�\ ��i3�|)sՀ���`����h��;�_);�ik���b�Bϱ�a(􆿳�ټ*w2�56kѶ���� �؇�M.98�{�����7s�9���o>��l%i�-5�e`��9�Zh|���!�`�(i37s�9���o>��l%i�-�u��Y'GF�O����!�`�(i37s�9���o>��l%i�-�����bp�%�)����!�`�(i37s�9���o>��l%i�-�����bp�@!�mg?!�`�(i37s�9���o>��l%i�-����n9�H\e1E��!�`�(i37s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7����n9일��Ѻ'N�c뵣�7s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7����n9읒��o�!�`�(i37s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7ݓ��E���p��b��L,d\P��7s�9���o��S8��<�J�QM�A�;�֋`N��7�j2�ٚC�M�����T�\ ������q�f@���#!f��O���H�"z�a<�Y�{'%s��.|Z���I7��-5��6��	���`y����@����gG�!��V�B����V+d�Z鎬������_�,��`&�;y!�d��Uт�d�٣���zR�K��I��� (�묈�϶�B��+ HY%T��BPAj&=�*$��
}oX�4(���k�G>Gqƶ*5�����e�`���;��|B�]�w\�O�bTG�N�����n��
/��y;��`2����]'\gWg��	�Z�kfc��2���8���+�^n=\f�5>���1ë�LA��R�ߋX8%�v&2\���F�`yx�>�+X�[�G���K!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2����97*�SCu̀A�pK7͍��|��W&":VA�ڦ�c4����g�Z��3��a���!@�f")z.��W�����F�P�7��S��h��d\�����l����� �'����u��r��;�jmT�#Q���V�_�mS8<�n�ݚ�Н��Կ���p5��6V�|/ ���we��0�U+�qbp@�!�`�(i3�����!�`�(i3����.��Ν�ʉ_��ݚ�Н��H����D�Xy����I/��\]� h�ҩ�!�`�(i3���ER�.0R��崰�7���ө�)�F��3A�)Oq�<sĐ!Eu��r��!�`�(i3p=�n��jP&}�m���V�)��>%���-ǫɒ�!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��Lt���hm�(��k8�ڶu�7�w�R���y�Z��T�.���j7��|�(�Zޙ��{�����!�`�(i3{Q_�dbzL���	%�3�
}oX�4(���k�G>Gqƶ*5�����e�`���;��|B���"�'Ŀ���Ӽ97*�SC�24����
�\!6�o8:4�I���c�90�Ǘa��xO.C�U��B��-��3�~\�0^˥�2����g^mb;�jmT�#bs��2[�a��o���zM#��m�!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}�p=�n��jP&}�mdN�<@Iv��nt=:�+�_0c ��k��^�1��dc�@c�����h�'�ɳ����Q�Y�;y��v��\���
^�ݚ�Н�:
��x�{�\��N�Ś�-����!�`�(i3�!AaiT��G��Hb� h�ҩ�X�o|3J;_Q���Qs��>H�,b�z'hۉ)��d�7�q�!�`�(i3����/uU!�`�(i3���Q�| EtT�K�b7!�`�(i3�Zj���
5/�V�q2P`��� Z�y��	����VPYu��r��!�`�(i3� �l	:�٭��W�!�`�(i3�̢k����^go���yGmϨ/��ww��	S.���:��-����!�`�(i3�Zj���
̲�2�!ڄ�]���J���S�<Ԣ�7Z�:1�\mdЧ^{�js)l໶�,!�`�(i3)P6����r"nCo��Y�d��n��S�<Ԣ�7Z�:1�\mdЧ^{�js)l໶�,!�`�(i3)P6����r"nCo[E�ގ-�k��S�<Ԣ�7Z�:1�\mdЧ^{�js)l໶�,!�`�(i3KP��(��6� ;h$	�kCF�(�����(�=�X���/��U�.P	HȆH�RtV�^!�`�(i397*�SCu̀A�p�����n���Ke��JW&�C��.��}Dq�f�!�`�(i3�5ߧE4��!�`�(i3�߆�p�h���/a�O<���H����@��	9צurT�B� �b��!�`�(i3�Կ���p5��6V�|��#������^�>������
�:qEp'{w#/ B!�`�(i3*�˜	����r"nCo��I�Ūe�ǩ"�4s2��ԜF��v��?���(�
nЯ�O�!�`�(i3H\wN+����&$?���I�Ūe�ǩ"�4s2��ԜF��v��?���(�
nЯ�O�!�`�(i3H\wN+���S=��-��I�Ūe�ǩ"�4s2��ԜF��v��?���(�
nЯ�O�!�`�(i3���v²*^�:�6�'�K1Y�q��؇�M.9j�֎���x��y�o�!�`�(i3!�`�(i3�����n�����h�&m����fJ�1D1�_'�脫:��
^��}Dq�f�!�`�(i3�5ߧE4��!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�3_�n^�	$m��M[K{ˉf�G�<��}�u�?�d���&��r
�ޮw��U�]��H��^�Zh$r�Eg�N>Zg���5φ��<�6�@a� ���N��ȥ�n4s1�U��B��-3��܌o�P)���L��mD���5]�7�癆cgQw�c4~Nr_�mS8<�n!�`�(i3!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"|�au�(Z�H<�2�8��C"���^E4+у��b�Bϱ�Җ���϶?� Zh�RG�p�P��c������>]&���F�x��&���ő��̼Y��7�:2��_
�u	{;jd�b:m�X`�7���ө$>��:</Sn��K��.1�e���b�|U�O�-F}���V6}l(f���r�r%)cA�$�+Ö��?� Zh�RG�p�P�"i<,��1��yM����Vm�:5A��p����E�El~pDa���UJaB�u"�����#�-�p�#8�"��!�`�(i3��ic)�̩*��c�d*qA����6\�4�@�� �-jېI�q������ л��E�BS�+��U�,�P!6���r����L�J)���� \L�1tSjv��H�������bO��M?��y�!�`�(i3��=m緒Sr��3��ő��̼��nF���<�W�.�P�	��
�Q�},\ͨ܉p�u-/���y�8��C"��|U�O�-F}���V6w��EO"�̞��>���I�Ūe��Z�Y� �ݚ�Н�[�t��#�Β �r��!�`�(i3�^E4+у��b�Bϱ���ԜF���v!��c���w�K����+��dЧ^{�j$��XCp=8�b(��Xo=��-K�!�`�(i3i���ؠ��6���9�
z�.�MJ�A7���ݚ�Н�t�R!ME�б �A	�!�`�(i3'�^�����ݚ�Н�.��fReU!�`�(i3�\d:0�g���C�U��.���|e"�� л���S�	RN&*�8#u���;�jmT�#��ݟ��Daa��o���T/Pr
�ҙ����l��.�B�;�ez8�US�B�!����r�7���өzW�&��F�u��r��!�`�(i3rI�F����ez8�US������`�K7͍��|��W&":�ݚ�Н��Ra])n#���r����!�`�(i3� ʋ�aGM�о٫��@�&����u-/���y�8��C"��6 y2��R�!�`�(i3�5ߧE4���ݚ�Н��H����� ʋ�aGM�о٫��x>O� &-���xԾ�J��RQH�RtV�^!�`�(i3�⵽2�RH<�2�8��C"���\hw�h��r�r%)cA/�r�]/2�ݚ�Н�!�`�(i3�#}�{�@�m�W#��H��dN�<@Iv��nt=:��:5A��p!�`�(i3��jVѭ@!�`�(i3�'��o�u:��_x�H_��#��SÚw�K���p��b���ez8�US�(_eW}D�!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě���ž_�FȪ���l��.�B�;�ez8�US�B�!����r�7���өzW�&��F�u��r��!�`�(i3��5��(���Z��oGM�о٫�Y�2]%�IG�p�P�m������� h�ҩ�!�`�(i3���(��K��.1�ޣHV�v&
`�|��K�z/�r�]/2�ݚ�Н�!�`�(i3[�t��#�Β �r��/ ���we��0�U+�qbp@�!�`�(i3!�`�(i3i���ؠ��6���9��,�tј�T�z�D�R!�`�(i3�	��x��ݚ�Н�!�`�(i3[�t��#�Β �r��x2%0�զ���Tٷ��1M�.(*��!�`�(i3!�`�(i3Y[�Yy�l�Y�F��(�}�1U��VP�h��;�(_eW}D�!�`�(i3!�`�(i3�5ߧE4���ݚ�Н�
�:qEp'{w#/ B!�`�(i3���Mڷ�2v.^࣡N���)x����J%g���ި���?�'���g�p����dЧ^{�jJ�lҾ�!�`�(i3$f��_Ub�F�S�1 �
�:qEp'{w#/ B!�`�(i3�⒍~����R��:�A���)x���3n����(��3A�)Oq<�WK�9!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j���_J��`L��Y-1ף�V�On��Vy��s�P)���L����
�\!6�o8:4�I���c�90�Ǘa��x���+�^n=\f�5>�gd�a�"�
R/�Ū�������f�YuA(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R��-�E��%�w�=�J�5n��>�my$�N��o�/���;���Ȋ�?Ӗ	W��e.�9��T�z�D�R�k'��e�ؕ�22�%��v�ک���@|����^a�nu4Bޗ��jw�	��!�`�(i3lG%��`��ǚ��ظ
��@�U#�s�Yls�<Ԍj��_�mS8<�n�ݚ�Н������y��'����u��r��`
 ֢���@�k��}!�`�(i3��nF���<�W�.�P�	��
�Q�}`
 ֢��.��� �Z��2S �J�A7���ݚ�Н��]��W���Sd�[��I����~u/��kOT�Ra])n#���r����;�E����T��O�T/K���r�����+��9,({~1JS�K{M?��y�!�`�(i3vx��c6���J���뫞ic)�̩�?D�8��!�`�(i35��
�4v�*�P��a\Y�����J��RQH�RtV�^!�`�(i3̲�2�!�����;q�{_8�Y��=�}�Vݨ��}Dq�f�՝� s�#���k$ !�`�(i3���D)��J�a$�Y F�*3��1�?�+��~!�`�(i3$f��_Ub�F�S�1 �����l���b�2D�]#�'"�8�5�� h�ҩ�!�`�(i3��|>�ğo���X�u"����!�`�(i3�߆�p�h��b�2D�]#����h�'T��x.�Knqd��^��R��ӟ-�%�ɍ��=!�`�(i3`
 ֢��.��� j�H]�����x���b�!�`�(i3h,ID��.2�6� ;h$	��*W�У�&-���x�'@�(��P�G�p�PXI����|�ݚ�Н���6����Αk�]I���,��~�\-{���!�`�(i3�k��^�1̲�2�!������ʟ��yM�B(p`D҉̖�7�j2����|��H�RtV�^!�`�(i3;+�'ն�%H=1b��?��^<�w�!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹��a#PMo�ez8�US�_A�IM���e���W�*�(4	d���U��)���Y;e�iKI/B޾Pb�i0[���S�J\7�_�Ƭ7~6O���N�_�ɬz!�xjzӝ���I(͂�'�ɳ��!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2�����G��!�`�(i3n��뾦��F{/�����,([�y�""p�2�ξ�b+}y[�k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}�:
��x�{�\��N�Ś�-����;�jmT�#Q���V�_�mS8<�n�ݚ�Н���s8��J�a$�Y ״$(�>g�!�`�(i3*��^�"~HR�3]� *�/��kOT�Ra])n#�V���p�H����<z'�$쾹KK���������E�El~pDap��k�Ԛ;+�'ն������|�Y[�Yy�l�Y�F��(�7 �E�!6\�
 �Q7��H_��#��`����W��yM� :H��\��v:�9
�F;p�	+��Q��:~�W�J��R��ӟ-�7l�A�A�dy�.�!p��q\sv�h��;�M)Z)�	�g ��-����!�`�(i3]a%ڔ�����;q�"��ӌ�r!�`�(i31���~!�`�(i3��JתMܥ�I����~u/��kOT
�:qEp�;�P�t�5!�`�(i3��$�B?��fg�p5��Q��"��h��;������Uxu��r��!�`�(i3�#�l+�����p�?D�8��՝� s�#���k$ ��'T���+��PJU����-a0a3����|e"fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�����REJm�Wd�<�g�DP�`�@s�U$��h̷_��yC��S8��ʹ}��S�٫E!��(���B���ި�����|`��'��>�4Nu{ᵿ���C?�Q䨈Tf�)rY�Ǿ{K���"��є�k�l�g7,I�@�"|_�8���< ����wWi:rö1M(7�������Xa������>�v�䩲$��8g�7L�k��.`L+�<f��J��׵�"0V�6�o8:4�I���c�90�Ǘa��x���+�^n=\f�5>����Db^5���0"O_�r$ɓǃl[�Ƶ��I�q����!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻt�{#	�x�H\e1E��J�a$�Y dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(�8�u?��I���?B��#Ɵe�*|�÷�Wе ;�jmT�#��"����G��Hb� h�ҩΏ��^Kho�7�j�Γ��-����!�`�(i3�I��m�]�{E��7ue��0�U+�qbp@�!�`�(i31���~����l�馍�!S��#o�]�ʄǡ��_qͧ!�S_��';��#j�ݚ�Н�?V��j�c�]���4��F�(=�ݚ�Н��̢k����w[��r^�.���ZL��-����!�`�(i32W���R0R�8�C�w~���Ѻ'yrf]���ቅ�%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��jCZ�zk��X\Y��k3�\��1A����>:��2�vφ��<�6�@a� ���N��ȥ�n4s1�U��B��-����A�;��27R���\���F�`yx�>�+X�[�G���K!�`�(i3!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}���=m緒�6�T5.Ze!�`�(i3x����E2b�z'hۉ)��d�7�q�hs�����F;p�	��Œ��S/ ���we��0�U+�qbp@�</Sn����+hX~!�`�(i3����;q��b+}y[�k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}�:
��x�{�\��N�Ś�-����;�jmT�#Q���V�_�mS8<�n�ݚ�Н�|�au�(ZԵD��0�rJ�a$�Y dN�<@Iv��nt=:��:5A��p��(1l�jG���Z��o�g� `�1KE�g�������(ӈ���m�r����/��@���@!�mg?!�`�(i3k���������|e"��w�w:�!�`�(i3��=m緒�6�T5.Ze����;q�#}�{��8y�R�Vyrf]����;�jmT�#��ݟ��Daa��o���H�RtV�^�'��o�u:��_x25���w̷_��yC��S8�~$�n�@�F;p�	+��Q��:~z#��#���%>�rGO�D mWN!�`�(i3/N2~-��x�f7﹏x2%0�զ�_*�`�	���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��jCZ�zk��X��%2�/�Cǫ��3ӀB��+ H� ��U�_:GK	/�en!�`�(i3��x���=�n���Q1���`����OP�˟<L�9�8꽻{Zٜ=bfL0S�t?�:��j�g�����_���Y�{'%s��F���\&.����ȕq��N�P��D�W ���!���c�A�L'�D�h�H�!yg'�UH "�r4[�H����Vhx���� �is@�����]��t�iZ]XF�hx��G��Zt%��m&<2O!j����x��B5�!�`�(i3!�`�(i3P*N�2���������,�ttT�r�pΚ�w]@� W|`f!�`�(i3�&8�,������k�v2<�����hWK{m35%,�!�H<�!�`�(i3�X;p`�V�׍A�f�?ǉ�=��<E�f��V�mK�b\��Mh�!�`�(i3�;�����^��&X!=��hy�/B/���^!l���Z1�:�,x�~!�`�(i3,54��]��)�4!�u3v��U�DnK�]_!C6%K�pıN�c뵣�&8�,���c��Vtk�)�p�X:��+�S�9;/���!�`�(i3!�`�(i3!�`�(i3��4MT2g��H#�"8��=�<���� z!�`�(i3!�`�(i3!�`�(i3X�PC!`�|��K�z�&�C�/���Y�l,�x�6�
X!�`�(i3!�`�(i3����+��c��+�y�^v%���z\�m���Iϕ������z_۬=�!�`�(i3�&8�,�w�Qt
����+g#>�����������622���k˗S�d�!�`�(i3!�`�(i3t<� ).�xz�\�{<S:H��+܆��K����!�`�(i3!�`�(i3-��<�ξ�\zǣ©���9��^K��[N���b�����sd�!�`�(i3���K�7��ãx���`</Sn����e���W�^�|n�M�!�`�(i3!�`�(i3P*N�2����������wbk�$+��m�yo���|��Mb��y9xO�`G��
���9	�Lģl屎�q�~�Y���(�}�Π�cC!�`�(i3!�`�(i3!�`�(i3��������+�y�^v%�������>[H����&?�!�`�(i3!�`�(i3�&8�,�-��A������t���hQ�GvE#�n�%)�ak�m6!�`�(i3!�`�(i3-��w¹��<d�,��L��~�Y���(��U��?D��!�`�(i3!�`�(i3!�`�(i3�F�7��Y�
�cc�V�/�"�����_G��?u:�L��!�`�(i3!�`�(i3w)����*�e S]#��+qѭ�+g[�,�ttT��������!�`�(i3!�`�(i3�&8�,�;�ږ�)kq�ށ �~����as��!�`�(i3!�`�(i3!�`�(i3�bV'�&�f�?ǉ�=����@!�`�(i3!�`�(i3!�`�(i3�U젩`#�4>?� �1�s�٩�����w0�!�`�(i3!�`�(i3-����b=�|�\m��l�eo�!�`�(i3!�`�(i3�&8�,�{Z�{0�;?7�k=��#SƏw0��;%.T-��!�`�(i3!�`�(i3!�`�(i3
�n��E3�0����</Sn���Ӎ�g�c�!�`�(i3!�`�(i3!�`�(i3o@
i��@f�?ǉ�=���P��!�`�(i3!�`�(i3!�`�(i3�����Jw����f�@�_&!�`�(i3!�`�(i3!�`�(i3-��o�]�S�*�K}��C��]1�
f5���lTN��I���q�}�('�Ŏ+k�n�U|��%w&͏��姸Kk	|���|<:����fS��j�ƥ��{K�	�~(�p��M�3e0�glƈ�|(G�$�E�#s���O%��>�6�t6b�x����7V��X�`�ƶ����"?��A$�P������5d��n4s1�U��B��-%G��^���x�}�yW���"sS<�0�zG��� ߛ��u�ź���4AL��άA�
����{_8�Y��=�}�Vݨ��}Dq�f�֌��-�a�ݘ<�̆xƍ2���l�[�ɝ���q00���龸b+}y[�k��^�1��dc�@c�����h��-�����s�Yls�<Ԍj��_�mS8<�n�ݚ�Н�:;P��� "���
w�j(���^:;P���^��w�����vo��Xl-�"���Yn���^S)t�  �@&�$���\��sȸ�"rR�H��c�L1���`����?��[��bq�q������Sz�����9�O��F���4AL��άA�
���'MtZ�R����Fz���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ&kT҉­B�0����3Ah	)ޟ-�b�+�