��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:��ښ�1oM�U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]���<�j�C��`��L&`^����8��U�Z봣��D��L���_�L�3��0I}.�ANMs����Ѡ�/�Ҷb��N�w	*D���y&�f��+K��[y��ڂj�x�z:I(wKq���/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�0k�5k��J�|(���u����l�|���j�I�?g�f��#��� �bRw�����IL�+�{Dr[��=�^S���Z���y�ۘ�G�|0$��&�^C����Jw�)��Pip<ɯ�nefR#O,.�c�u��QF}����;�A3�'���/�k��±'�R��;L$]��]{�[N�4�=,����Ϙ�Ԕ'�Ӝ[Y NoC��c�S+d?S�7�$�>Y9w0�R<�CW���V��r:O!�`�(i3�g���}���������8*��#�N��O���:�9`�p�0��&�����¶	�Ev!�`�(i3!�`�(i3��1�<����>l�ݯ���9��)����6q����"� _�i��i���5���6*�t��L�kjt���?�����Jm�W���K���v�7��٤cF�Vq	�!�`�(i3!�`�(i37p�J��PW���3���D���o�i2��0�ּ���)��G�������ϲ���>h�c}����>I	���(��B�:����@���4W�-c8��"�a�O>*�ׇӭ��!�`�(i3!�`�(i30R��=	�@����W��nl@O4茸z���q����R��C���CS�� ��!�`�(i3!�`�(i3�0�9&،EB����n��|1�b�YL��&\VI`,xJ�����gc �{�=2���p�)U!�`�(i3!�`�(i3X�o|3����x�u��"��휺�&\VI`, �DO'�L5я�����0��zO�)v��$�Pr`7ï&��.�-�&��4�%�@V����S�����Ŀ"���J���>�$!�`�(i3!�`�(i3H������gf���5��x��X�mϒ����y��f������E\/P*i��!�`�(i3!�`�(i3!�`�(i3 ?[n�:#G� �b�H~V�I>1͊���3-���I T�+����̵��8<=!�`�(i3!�`�(i3!�`�(i3C �@nk�@���;)�����<j���ֵ�Ů�y��ͮ5��}��6�8�-Zy?X�`:;��
c��@*1�L� ;N>�G�$U��ިB�Y�5J��5:5J��(�ߜ1�ׇӭ��!�`�(i3!�`�(i3!�`�(i32g���`����&\VI`,J����^��f�������W�� �!�`�(i3!�`�(i3&��潹��a}	/ȸG�$U���pJ`��8������O�w�V
�1!�`�(i3!�`�(i3!�`�(i3�I��(,�a]�l4���?�AO�]X��ƞ2�� u8�"�6���G��ꚕ�(q!�`�(i3!�`�(i3�EH�2�L@���_r�Gl��c��#
Q�����zwK35���h�w�)ꣴ?���X�!JFh�`������eC����	F�o�=��KQb�KK�y؄@�!�`�(i3!�`�(i3`RXK:�w� 1ܮ��gf����;��@B�a����K/tE@��j�g��o��,�r8ЧڜX��hvծަ� �0���o���Ѯd.�6��S�6�0RD��}��b.զjUǡ�9�ă@���3)ͰnL
sȸ�"rR!�`�(i3!�`�(i3�z�:>�=��9�V��r�-b0��[��u�j��-xIYBN~x~,[ӝ60��,o�!�`�(i3!�`�(i3!�`�(i3Eu^Q��X�[�"�k�fQ�����z�xO��̋z�:pF��w�=���6�t�qŻ
p�!�`�(i3!�`�(i3!�`�(i3k��U_���nཱ�&������!�؟�r�Y�}94�h	U����f�7U�i�#!����P�>+�va��2	p���>/:ܝ	�@�ׇӭ��!�`�(i3!�`�(i3�>L���L�ɚ5���x�[�%���%���=���pw�ۢ2��vR�J���}���	��!�`�(i3!�`�(i3����N����������(��K.���ccnh?��7>�����D/͘B���&,��*eM�����3�j��~[�h��\�ڰ���gLE�z�K�y؄@�!�`�(i3!�`�(i3�>?v��B{?a� ~>J*�ya(�$>&�.Q%�i
u����-1<@GŚ�ׇӭ��!�`�(i3!�`�(i3eI �#��I_h�R$:7��}�؝�T�D24N<I8����\.Wֵ*&E�^8��xt��:_/�~8����A�߲wLB�w���#✲�@�킍�"�?���Fz�!�`�(i3!�`�(i3�s�cn0�u�A�qL��D24N<I8����\.W~C*B Ɣ��(J�fŊJgSᚄ�j
��a��ǂK�O)��+`�{�gt�R2���4eM����;�0Z�8��1	/��R2ռ~�S�N�\�:����{����~��➛����Xw�e60���Ϧ�lـ��Z�>�=��$��6��{ֱ@���O���:R� -�*3fх�-�@���q�qp�HTEn����1��7��w׸[�	�+%�����;�e >�#�mi��,�kL���Pv�����'Q�@RͤUʐ�{?a� ~>�8�<��{�#:B�6��1��h浏��������S����3|��@$�g�9f�oF�7�8��i�c�������7>�����D/͘B��)gI�qd��+L{��+x⣗�C�|�6G�"	�WJ�Slm���`�7^�	���*�C ��s�Ε?�������4��A�Ww�=�d2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hͥ<#���vSB��n
HDW�Gj��o�/��];Lth� �K��G������\ͬ�W����]��Q��S
�yl}Vİ�M�W9�f^�Ԫ^��rL���	��D9�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc	���[�;�4A�B�'���W����+n2Xh?J�k;��7
��t^�L3��헙��l���Cf�O�P,&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q��f�SR�v�����������\͜��ͱ�5�����\�� �K��G������\����h:�Ê�����\�$90�H1�����\�P��y40�^�����\�T��v�`2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������w'��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:��ښ�1oM�U���T�����\�4�s.)s:^�e��Vu�?*t�ML�#
ơ)Ճ�v!�zg�Z�$�0�iH��V_@mv����`K+b�ĈPR���"�D�u���ӹ`^?�rfS+���RL�a)	�n-�~F�~篟|�!?!�{><9�U���Tџ�_�v%�I �"혱
>2�%1[br�O��C��0������m�Q�pY�� e���T������w�>��S9�����}ZFȑ�R��>=�6�'�al��p;��|B�\,הE�_l~�[�'��l��Ҥ��5,M���p����%����L9�R���\�4�sp�3��I�BK9�H���V����U�[+jm��Sd,�ϱ�E����}�?=����u��w)�S-!������~篟|��*�A���I�n����fџ�_�v%�~G�6֍�r`_��*�u��.t�5�M�1�>�8B���<{��*b.[P�x��t*�=�V��u�/��m��@��V��=B��,����t_Ȥ�W�w��fD ��b�FP& ?[n�:#G(+F�	BaN恔� 90'�f����&�&�
.�n��������SiC���\#�t�����ڕ�>���??[�o��RL�a)'r�Ӟh� mߍu�M9�ߤ����Q���@m��7C��H!�������0�'+��h��=o����"���	x]�"�PL�,eHc�J�M=���-�:1,ĠԜџ�_�v%�_ y�+�3F��m1G:��"w[&�K!�#n��]t�#K�{�:H7ǫ�V���V�/)�Myիnň��h���|~�@����k�8���҆�|n��)8P�d'�%��hݜ�����AQ6|U��<d�L\�Յ�B�U�٣�R��$���"HX��+��^gg1�
հ��C��iF&�A��h������:��KL�����.jB��@۩�����k�8���҆�|n���&�]�68��hݜ��  Y0�����N��%L\�Յ�B�U�٣�R��$���"HX��+��^gg1�
հ��C��iF&�A��h������:��KL�����.jB��@۩�����k�8���҆�|n���h��C d��hݜ�����aj)�>�,r�F@�4%������I�Z�*�I���Ϊz�&���Ḱ��fM���v#n�0؈sU����A����&D��0H����RL�a)ѻtUWR���I����gy3�]	��>	|!�zg�Z�$m�a�gPM��r9t���k�8���҆�|n����{y�ڗ�B�����[AF��ѕ���<l���9��Q��CpC���D�v�{���c�5��<�>�N��̴�*V��z,L���	x]̍��;������#x��(��[�� +u��Ix���y+�����S��&h���y���La��;���g�Ȝ��@�r�O��C��0��$�>��w�*��D����Ǳ����w�>��SX`X�B%�r���7ȓC�-`�e�g��!��x���� �"!B�������.�-���
E�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�f<�,=K�F�~�����J&���f<�,=K�F~�?|�[_�qR!��HΜ._^���^��bg~/�ח۲�J�[j�fTܷ��WL�C�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��P��'�<	�\�Z�م2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR@�/-��E]o��in�m��+�<4��ˌ�ň��h��j�V��v�����>�Rh�&�~��e hI�ˋ��vE-,b����Ǘ�Y!�`�(i3x�]�V��ι��QG���/�}���1�1�ҕ ���3�ҺIÙ=�HF���m¡Cd�_���+��;"�g�E����F�'n�^0o���˟y��)��'��8�-Zy?X�!�`�(i3JHn��z�/ue:�<� �vBX�y�`4Zp��/�����Q�^�y�zL͊�q���Vǃ���*L�E�w�̙	,N�����JHn��z�w٩L7��HUv�׿e_=����Y.�J�4�e�(�4q���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3����j������)���g�{V�b!��u�$M�Q���?���\z-����o���������i�A( ����_ֲ��mŹ�[�g�DPp��&\VI`,�=JK�t0�`v!�����h��*��{m��=��9౲��+�J�������V����(��ؽ7$�	�s}��[	L'J����Rb��Y�W,�KYeu�BY{Y����H���/���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3i�/�
���)�����`�-�q�/��s'�\P�����i�X!�!D��(J�fŌ��P��\�v���GAџV������!���C�/�yT��H����7�ܥ��2��t��m0����r'��˝Sz��E�4.@��n̈́�zL͊�q���1m��d+0�l�R<�q��f�}��h�'f R�E����F��j��\w��0]��0�&�ͭ�h�O�0c��Et��q���U�C#/<���q�VP��@�����ɧ�J�8�J��	��	Mk�rN�By3��<�]�!����M[��Ǣ��aX� �䓒��x�O�,�j����0��G�4?�@IE�U��>��l%i�-�%t̓�@���I��gs7��-��%Mό���.Ӂ��̰�!u`Ʒ%k�����
L'���Xw��E�d��7#1=��*Yl���#�]�!����M[��Ǣ�7�]X]��@��$�K@IE�U����S8���IO,�?9Pjp��}%����͋�7>�����ǚr��y���Δ��p�T�\ ��֕ߝԀ�ح8Y��fU�aB���$�O��1���H���;��"B��$I��w��,c�A�L'Qī�*pY��am��	t���o����s����|#9��Ė�{�!�`�(i3��(�
t�������2%=dϖ�i�q㧵�0������0��D��L���_�L�3��0I}.�ANMs����.S݃�0G+2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Pc,�w�&���#tvQ2�����\�w�Y��k��ı���$��������j��t�w�c���������@VF�}�
�?����Y�l,΁�a�n��JHn��z���i{8�.Pl�:����Y����F��%Ah�%4
>��`���oHe�-�c�n�c��	n�E����F�_���˸@����gG�v!K��>�Q\�p7s�9���o��S8��<�J�QM����2�E~�����R��v	�R�wX��}�
�?��(R\֎u�eK�	�$V��d�٣���N N�S���c��:KY7#1=��*��i%Q,$'���Xw���,D�H�p0���5irAz.l�n`5�fK�\w��0]b!��u�V@���gx2"�,�>E���]�!����w�Հ�$����Sr]�+^g���+�J���q���U���g�,P�nw�����A�?���0yV�6IWJE�!r}<ﷹ�t�Z�f����@1��?�T�\ �ͻIb����rs�i�/ �m^'��D24N<I8����\.W^�V]��}R�wX��}�
�?�套�qD0t
�X��)�Bh����YW��b'�3Ai�@����gGp�E�H�+�(�9(��Z鎬����z�֐��D�iI9�o�L~΄gO�3��|��[��5��S	JZu`Ʒ%k���}o�@EZ������i��.����.��$�\1^O��[�~�����\1^O�Y\a�A�����d֕%t̓�@�ۅ����*���n,�d�5)��Z^��i��.�w���H���;�(̚N�:R��1ig!
,=����I�1(,.��FҼ�^I�R'cf��i�X!�!D��(J�f�w]�IB[�)����]�5�O�%E#P�%t̓�@����Edb��7>�����ǚr��y�_��wBW��y��e��#E��δ�p��������s��� ,��rQPQ%cp��g���t�]V��	��y ��f"�7�]X]�O���&��G�!���(�Ea�7�φ��<�6��ً��:+"0H�=ϑ�φ��<�6�V�ҁGGSoJ̈��:��:���
W�&��9Ԍ�����!�`�(i3$H#Ö�U���KX}�!���ra�[�k(���"H�@�өN}�m��{W`�v�L���f70���Y%T��BP	�I]����2N��n�F���0'��=���ł�"�,�>E���]�!��	Ǹ�y85�C��H����Q^�MY:�6���;b��g��U-�e�,���6+� ��b�FP&p�]f�"v!�`�(i3�5c�;�K ���l�;���EWr���gRI/�f70���,ԯ���gnņ��#�b��~�26��\��`t�B<4a@r�b����+�J����uݯu_t����Uh1�yO�E���%�;���EWr���z�щm�����?A����cfoa(􆿳����{��~�26��\E;�����!�`�(i3X2zӼ<�z7�g�+���ֹ�͈����$�Qu��`2|`Kr�|�KT��E����F��Op�ե[��GAџV��$�Qu��`2|`Kr����ڽ0��E����F��Op�ե[�u�,�sޤ�$�Qu�ْI�s��N��}���:�Z�{^}�=Ll���Pʶ=��݉�h�B��.��|ȃ����qD��=a�^7�1tSjv����"sS<6Z�٬�[���e둼�;��N�����1tSjv�.��J��X, ؖz���q9+t�}�ݚ�Н���$"'�ь%�"�Z1�j�,��f;I"����5'�wbk�$T��8$2OU�1Q�\��^����!�`�(i3~�`cC�4��5��R��/
�zS��j������!���}Dq�f��?�_�+��%�"�Z1��2�A�dv9�]�REu��r��y��j��k
�X�nZ�l^@ !M��SJc�=Z��}Dq�f��� л�V��w�G��S&ϊ*7�xs���ݚ�Н�����a�~9��tf��!���gRI/
�T�r�5�9��n�7�Y���X�q]���]�o��Tg�
�:qEp'{w#/ B<�6�Q=۸v��I�TNr8�ȭ�z¬��p�m����ۗ!�`�(i3�S�Ĕ�ZӇ�;tY���?EzIA�M�d?�qo<�kh>� F��9�{d������Ө#��^x�E����J�UE�lN��]۔2�/��@�����%~��bSo�3=����|e"�=�<��=��?����\��;�,���y��lD�0�+i)���{ֱ@�G�>�o�5�)����k��O4��ge5�||:�-4-�9�����T��� �bհa%�z���vo��-R$��{1?�a�uE9�+�����vo�H�-��
�$��^)B��B�嵧ܵ����s���<]���}Dq�f���Ě�����}Dq�f��5ߧE4���2��}��E2�DZ�⦫/���bxK7͍��wAA�Ɓ=<�W�.�P�H,0pMp!(@X~�H:��1�, �����{���}Dq�f�=�B4˖�J�a$�Y )P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^����S`t�L?t����}>�O���(%�Υf/�|�R4�(�q�N�ǽ��B� �b��!�`�(i3O���8z����( k��o�{��Ļ�*�@;��-b�uE9�+��;�jmT�#��'}HڨF�:v�ֶ�����Qi�d����VZ��1����C����"� _��J�8^��u��r��!�`�(i3XIN����w���B}�����z��](g���М��^������*9�hY�%Ͻ�w���B}0/0`9N1�B� �b��!�`�(i3�H�����7>�����D/͘B��< �b�V0e�{�W!�`�(i39�O��F�`,9�H�W�I,�D�y:#9�]�B�_��wBW�MM
��,=*A&-�Ri!�`�(i3�/��@����}���r$��^)B���)/��:5A��p!�`�(i3�H����-tG�r�Β򨞊i�����-����!�`�(i3!�`�(i3�q�	��c�/f���H�pG�}#Ƿ?j^y6^�!�`�(i3!�`�(i3���/����n�@�N�m�[�N�:5A��p!�`�(i3�wӨj]h�O�M:R	� �}�휨㇟�})�1�Ʉ*R��!�`�(i3
�:qEp'{w#/ B!�`�(i3�y��j��k
�X�nZ��3��%�
�T�r�5�!�`�(i3�wӨj]h�O�M:R	� �}�휨�]�!��	Ǹ�y85����[����:�[�LH`y
��1��� ����P�7� �:5A��p!�`�(i3fĉ>99��A0ok��!�`�(i3���y��lD�[�D���ϴb��������r-�P�)������юw᥽ ~뀇ϡX��:���P�ݚ�Н�!�`�(i3�g�`2|W	"E&��� ���������t7b)J���9��V�9!�`�(i3\���F�`y���%~���^�u5��-����!�`�(i3!�`�(i3Z���ֳ���Zv���;��K�p�9"I�����眯}Dq�f�!�`�(i3HN��R��bP�63Z�t!�`�(i3HN��R���מu��� �H�0��
!�`�(i3�����!�`�(i3�/��@����}���r$��^)B���)/��:5A��p!�`�(i3��=�g�żפ	�?9Pjp������PN��7�v�ԯA��bu�x��ݚ�Н�!�`�(i3��)�hV�|��L���ʭB�?�`u��r��!�`�(i3!�`�(i3=aUh������zbG�ZVٲ���<���!�`�(i3y-�S��E��*��Sx֐�M�4m�ˈk��Z��ݚ�Н�!�`�(i3?V��j�c1����?���L)��{TN��U���'��L�xt!�`�(i3�Ra])n#���r����!�`�(i3�wbk�$����$��s��K����:5A��p!�`�(i3?V��j�c1����?��&tS�D�'���Xw�j�7��Z�qҪc��(jy9d$���?�y�B���0�&�����ݚ�Н�!�`�(i3$f��_Ub�F�S�1 �!�`�(i3�H�����8�ܩ�òo�����=������&G!�`�(i3!�`�(i3�<�W����6	D�NQ�4Ư�ƧE�f�s�#>������!�`�(i3fĉ>99��A0ok��!�`�(i3HN��R���מu��� �H�0��
!�`�(i3��Ě�����}Dq�f�!�`�(i3����0��Gd�~{��״$(�>g�!�`�(i3$f��_Ub�F�S�1 ��Ra])n#���r����<�6�Q=NUl��F���h��t���>������k$ ����l��	ͰZ����XW�G�<I�^$D����(R\֎u�eK�	�$V�G��Hb� h�ҩ�!�`�(i3�(R\֎u�eK�	�$V�n��뾦�!�`�(i3�2��}��E2�DZ�⦫/���bx:�HCaIMl�mזc�S�!�`�(i3��jVѭ@!�`�(i3���̰�!w���B}�#QSU:�����|e"!�`�(i3套�qD0t
�X��)���nF���ܙ�[-<�+�my$�N��YͲ�!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN՝� s�#���k$ �� л�����W�bհa%�z;�jmT�#�G�2ޟ'�XW�G�<b~*��s��(R\֎u�eK�	�$V��eu�j�~�e������5)��Z^�d9=���u��r��!�`�(i3=�B4˖�J�a$�Y ״$(�>g�!�`�(i3(@X~�H:��1�, �����{���}Dq�f��2��}��E2�DZ�⦫/���bxK7͍��wAA�Ɓ=<�W�.�P�H,0pMp!
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�g��ޏ�Jw�)���%������`u:�Q>�5�Y�w���ؤƂ��l�O�{ Z)*Q�]�(���V8zA�k��~��/6�o8:4�I���c�90Mj�dL�{y����i�q,?5q�0��g�~�
��lnw*�r$ɓǉ�.y�U=������&Gџ�3~�l"+�B-�D^օ?D^���k��^�1��dc�@c�����h��-�����s�Yls�<Ԍj��_�mS8<�n�ݚ�Н���B/�w���B}�����z��](g���М��^���'ƃ�3�Y1tSjv�����l��i�	-_�ވ��*I���b�Bϱ�}���yb���?\MP!� u��r��!�`�(i3��V8zA��ִ���	��ݚ�Н���w�w:�!�`�(i3Sƽ������B�% ��g3�q?-O딈pᜯ}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}�7���=�X�
j$�h\K�5~�������g\�u��.t���r�}�.��1:�p����ǽX�,4�?nϦE�6���Y�`(ggE��(G0��:Ȭ<?L	�φ��<�6�@a� ����C�'�ą�n��N��&jc :L�j�N�zg$]��0�N}�m��{W`�v�L�Ⱦ������<3C���_����$�Qu�)�˥D@��'T����:i.ߋg���~�26��\�v�F#�5�#��P`����KB�c
5Xn�DIc�&5�/hy�b�G2��$�Qu�F��&��1�����Q�X��ZG>�A�/�����%>%�����+�^n=\f�5>��q����.ǈ�����2G�,��R(�U���e��d9=���u��r��8��Aꗇ���@z\��}Dq�f��o�D:dǊ�� �������#M&1I,��,�\z��V��i%Y��'��_�]��_��0kB�����Xpn��2J�cFQ+��1%��*ȑs��-�������vo�H�-��
���Ӓ�ap������T냤�ME@��j�g��o���^ԟ2t�VݝH�2d��ݚ�Н������]����o7��	ڊ��
��
��zq>�ݚ�Н��� �?CtY��zek�GHn�2�/Xw�e60�W��[8$h��/z_�����h�[`���|C������f_�������B�Ra])n#���r����Z��JP��ꉂ��dC�؞�W�}U~܎VV��fĉ>99��A0ok��$f��_Ub��7��G_��k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-����;�jmT�#�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<b~*��s�?�����&*rB�WD�{͘6��q����1ig!Ir��͕� h�ҩ�����}����o�6����T٦�͒))X!�>P�ݚ�Н��V��i%Y��'��_�]��_��0��5�\"^�� h�ҩΗ/��@�����چ��N��Ưb75���J>n� ��V��G��<��
�:5A��p��6������S>��.��cZ���+���L>!�`�(i3���F1��kټ�b�	�RCJ�����@�ĵm�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�q����.ǈ��������Ύ�B$K1��ҔWohWt�_a��O)%�����r��y2Q�@2�C+��!��ͳ��[X��:''�$i��C��g:+�+x⣗�C��ҷ�㗼H�Cͩ����;nrZw�Y���q&A�Y�$����9�/����tl�d��/r+���Ã��\��q��~�26��\E;�����"�,�>E��0ϥ�IwYn������pV��+x�r�s�*�I�%.)�VÛ��d�������|���bF����~�26��\�C�LsM~�?A���"5� �Sd�Q�%�2N��n����:�j�������5������-"{b���~�26��\;��B�lX�i�+�ؼ�\�v��8&���I��S�J\7 ��>�:�e�;ed ̅��Ȝx�5W ��̫(� h�ҩ�:�6%��"��Ս�+Yٓ7���($�3��0��fD��j���һ��q0��Va�ir����0��G���_��b~*��s��(R\֎u��Gj7�uz-Ǆu
N��!�`�(i3�~m��p!)D�Мf������0��G���_��g4��Q1�BC���U�
{�~jYw߿���̙	,N��Y��)��!�`�(i3z�wΙ#C&U�)j�S!�`�(i3
_g��c��v������܅�E!�`�(i3U����ޚ�^�OG(�((�]�!��	Ǹ�y85��8��,	ij�i�+-������]@��2�K�,>0���0��Jn��ݚ�Н�m�ڨ�hծ!�`�(i34f��L�I��~�Tz!�`�(i3���ڍP[����!k��e!�`�(i3d0?�s]�[�oY�ՙ��~d�[��$�-�s���o�!�`�(i3%�yLp�h�C��_U]����9�s0��i?*B^`ٌ��(�ґ��:�!�`�(i3��Q�Y�l0}q{���}m �"�KY`��o�,�����`!�`�(i3��N�T?wZP���m̞��>�rS�b�8Z�����È���}Dq�f�H�����?�@,��V�ݨ.�ϟ�v� (��F�z�8#��v�9��!�`�(i3�N��[r�+x⣗�C���ё�^��� 7��{���������m��vn6g��El��.� n$fK�B���!�`�(i3>�WS�2v���� ;�ǆ�A��Tk�p�e!�`�(i3s`<ܧ��(7z����`4Zp��/4Xf��GH�RtV�^!�`�(i3}���yb��rO��E#����o�����[��l_!�`�(i3�5ߧE4��!�`�(i3��#�a�Ą���u�h1���_�M8���%~��#�8�C�	��-����!�`�(i3D��ng�.��5,M��Z&�ā����Hɓ�����f�
i�c�r�!�`�(i3�Hx&6��ѥh���>�
�E�6�g�Z~~���<�:5A��p!�`�(i3Qi�d�� �"7ۏ�+�-�����:5A��p!�`�(i3D����pG+�X.6���&��-����!�`�(i3<�6�Q=�=#+�
�e]34}�ݚ�Н�!�`�(i3`H��N�:�j����*;b�PiU���ڑ�H�RtV�^!�`�(i3����$�����F�z�8#s��qO���������6/��g7��ݚ�Н�!�`�(i3Z��JP���K���&��|��Ǎ�/(�1��!�`�(i3!�`�(i3���F��O��ݚ�Н�!�`�(i3���F��O��ݚ�Н�
�:qEp�;�P�t�5!�`�(i3Z��JP�����>�Q��!���c�A�L'W»��`�{͘6��q����F�z�8#3�N���[��}A?���`ޘr��!�`�(i3�k��^�1���gRI/
�����Z\�>�RJ�B�%3�Y]�|�$�������ݚ�Н��0�9&،��1ig!&k@C�Ɨ0z�cULE��K3�jAԢ�a\�%o�P��(�cR "�=���y�pkv|p!�`�(i3�y��j��kb��4��;J�[��?�8=�V�����������|HY�5Zє���WBe�������R+��*;b�Pi��}Dq�f�՝� s�#���k$ !�`�(i3�	y�z��k�)��qUv �6U�E��;�$�	�y�o�	!�`�(i3Z��JP�����rc���9*�g�ںOo��[*�e��,�g�čVU���ݚ�Н��0�9&،��1ig!׾ŞWsuz'���Xw�j�7�����P�|T�O�޿M��}
Ĭ��S��1ig!�l�-��;�:5A��p!�`�(i3�S�Ĕ�Z���d� |�yԥ�����v(*��娥|XK�e�BLL��fL�D��7C.9�����b��n���S�P��~�]��%E�!�`�(i3$f��_Ub����pT�!�`�(i3-I�!A(��K��ٳ�!�`�(i3n����Z # ?[n�:#G=ac9zAuHi�s>G!�`�(i3���'��@�my$�N���ڦ`�C>
�:qEp�Q�������;b�-�2��;�P�t�5m�ڨ�hծ��Ě���<F� ���Ք׹���C���N S������Q>��	�=5��f-�*��	1g��`	E؈sU����A����&T'	�eݷ�����k�ʇ8[�r�u��� t�Y@�Bo0F�Xt���#��V.9	sa$f�6�v��N���v|hsm�N�_s�=_xغ�#��@����T���Ӫ!�J��:����p�m~|���\f�����珶��JHn��z�"�u^��اHfCf��qy炍&5 �Q�d�l��5�9�=˳�m�
|�NwWkp>��C=��ʢ����~��th����ꠂﺯ����m���8�'\0�g�;�1Ȧ�8�'\0��a��i(}�
�?�4F�M7�ũ�}������Xc��1?�mm:��n4s1�V��o5]�|����qtM�,!h���gmJ/��{y����i�q,?5q�?|䞯H+;��.Ҭ�{�6�C������n/jF�ཕu�/��kOT �ԣ�e�����W�lX�,4�?nϦE�6���8"��l��C��MbI�)��Rd!rf�.Ur�����5B�ò+o¤�l���d��R���"�Q> ���8�_�6�)�E3	�t*�O�kZZ��&\VI`,�R��a[��K�=T�K�ꬠ$��0�l��o�s�"7��̳�u���4���?Q���&i����I�4Ca�6��3�����kN�]��1ކ6��3��%�~n0O�0��ݰu��"o�����q�5�p�mҷ}["��4��z��0���7z.��U���7��C�������i4뱙±#W瀁<�6�Q=E���M�n�� �1 l��5,M���ϸ����#�Tޞ�j���-�	B(�	<��	gv�\�˞N��� p{%AN[..�������z�U�n�;��sM������o�4��f�ŮT�*�ӂ�@�{�6�C������n/��V8zA�o��<���� ��V��G��<��
��)����y�(R\֎u�eK�	�$V�#o�]�ʄ�;4�zu%��XW�G�<b~*��s�F�KD�Vr[/}>5��0+�_0c ���x���
IyhG+_?wʊ��F:&�2�����ݷ�pB�ae ��[�S"�~L7T�s��R7��
�Ͳ��.罤�*�����:�I���Oj�\Ʊ��������"9V*K����0��G���_��b~*��s��(R\֎u��Gj7�uz�Va�ir��dc�@c�����hž_�FȚ���@@TN"����"�)O��ւ�Ѓ0�&�2�����ݷ�pB�atG��7��V^g�)�.��~L7T�s��R7��
�Ͳ��.罤�*�����:�I���Oj�\Ʊ��������"9V*K����0��G���_��b~*��s��(R\֎u��Gj7�uz�Va�ir��dc�@c�����hž_�FȚ���@@T�7B(�!��)O��ւ�Ѓ0�&�2�����ݷ�pB�atG��7��V^g�)�.��~L7T�s��R7��
�Ͳ��.罤�*�����:�I���Oj�\Ʊ��������"9V*K����0��G���_��b~*��s��(R\֎u��Gj7�uz�Va�ir��dc�@c�����h�E�i�m}6߸��S�Ȍ�?|䞯H���~�L��i^��quA0�e�?�Vx�B{cӏ��C|�����f�q4򿠺{��������y�:Fa�7������A�������a�(@X~�H:5irAz.l%��v����l�^!7#1=��*�#QSU:�����|e"%��7uJ�*��gB�����X�^>�ݓ�W�����zc�1Tٗ��
QV�H������V8zA�o��<���� ��V��G��<��
�-�ྜྷ��H�RtV�^���̰�!`�����'�^�����ݚ�Н����F��O�VA�ڦ�c4��
�`ja��1a^��ݚ�Н� Ӄ�&��P �h7D�v��ONH!�`�(i3�%t̓�@���ʳ�(�״$(�>g�
�:qEp:䩒=]'!�`�(i3�h�͍��&��8�'\0�䕀��jul����l��i�	-_�����>w��-����!�`�(i3�K�&�a�W�^�|�����NM���fĉ>99��A0ok���H������V8zA�o��<���� ��V��G��<��
���ʙz�PH�RtV�^���̰�!`�����'�^�����ݚ�Н����F��O�VA�ڦ�c4�-C��k�@���SxF���gg�#[�ݚ�Н� Ӄ�&��P �h7DP"G�wk���U.+"b4��ϗ�\�8{]dP �h7D�v��ONH!�`�(i3�%t̓�@���ʳ�(�״$(�>g�
�:qEp�;�P�t�5����l��i�	-_�ވ��*I���b�Bϱ�}���yb���?\MP!� u��r����l�^!7#1=��*���d�L����|e"$f��_Ub����pT�G�&ց�*�&��j���3��Y$�(@X~�H:5irAz.l%��v��!�`�(i3=�?��3�W�^�|��/��kOTm�ڨ�hծHN��R���
�Ŏ��Fr��j�W����P�k�P}ъ-���/��/z*q+6j�"Hs�2�	�L]s��ǿL��(���ћLo�"���8�ldF�$��A@�r$��^��
3~��+��Փ2��I��N�m��A�x^V�����b�| �t�q��?K��W�u�#!��׏��Z�ׁ��̰�!@EZ�����h��N�M���TB$�V+�B-�Dא �k/�ݚ�Н�!�`�(i3��7I��٪�E�d��7#1=��*���d�L��E�u�N���*�����:�I���Oj�\Ʊ��������`����ݚ�Н�!�`�(i3��7I���aT��3G?�d���&��]y�Q�'f�c&�:�ܦ��80	4T������'��7�@�0��:ށ�b��� ���풲m���<x!�g<*0�ݵd����5/:�� �L����M�,!hޖ�A$�P��O�@יߌ��omq��.��|ȃ����qD��=a�^7�1tSjv�t�R!ME�'�^��������@|����^a�nu4Bޗ��jw�	���|#HK���	ͰZ����5)��Z^�'����u��r��N
�����"ª�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��N��)��,Ƌ��Qk���l<^���H> �wt���+��\��y�`��vN;��Cٯu)����bX�d��-��!$
�d�u̀A�pd{��8ѭ���'xTNr8�ȭ�Vx�U�4�7�K�ŠX, ؖz��wl53�e�'{w#/ B!�`�(i3�H&&����Iihs[S@�b�F1Q+����$��r����!�`�(i3�p$Fi
m/4@�s Oag��.M=��<�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h-�b�+�