��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S���7a�k��rD?=N��J��S������!P7TǱ�J���G>[�{����iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lV�t�[;�Z��4d���Ġ���딣0&_���X0���2|	p��rw@	@us����p��Y?	��u|��yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��I��Sf	��,h;2���۟�
$�e
�9��Ax!P����9SA���S�BgV�0�ם�kAR�o	%1 T�V	�tL��	�<�A�}Q@���rah���"��yQ����D�z05��ϽE9�v'�P*܉�a	p�����i���@��a����|�9g$v.E�F����K)�'�K������u�[�ү�jcw~e�k�jz�����[�A��ǡ1M-!��*�;��[g����<��m@�k����8��0jx�9��	���9~����B������UE7�F~� ٦i�� <;y�r� ���InV�	��Wf'�j�"���M�	4��|A�U�O�|�ҷY�
0���ۭ�(��]�q���J�	���<�:�g�q�hu��m9g��گÉ��`��Cm{39��ꎸ%I6��_F19����x�<ttC�\�"k�-1��	-#�ש_P��r�I��T\��2ei�P�?���k��	n�#V�&�tٙ̃����
�t��b�`J�ǔ�Ɔ]hF�:��84C��i���F6����L����_ 7�̯��n�b[�B@|���!�:&	��/v�n�NQa"_x����ќ� =*$�+�9?�\�N̤뢲�
�v�����M	F���w?����^6.������aVA�J����,[$�
e{pY�w	����he,OL��nZ���g������
�lg!���[��[��尿��Z���ᡔ����¬W
�h��%��F�k� c��(�U�4�����j�|�9�������7fiͱ
��K��w�\��~����p�H�^⽂=#fl��@7s��f@�A�m|�Gw[	zF�N�>)c��Ѿ��/@���E�V�^�*��\0��L�P�XR�؈Ϗ�g8L���7iZ�]�å	��eeՂ�v3Y��P4n@�W�a�h�w?����O�"�F�g[�;�X\�Tpf�\0b�VQ��� Ua�,�	�[�1�"�k:]��9��4��ěyp��Ǩ�,�g�N=��Ѿ(G ���lXc�����/�l�{x=y��KO���LTɓ<�[//Vq��._�3�?�oxurD5�azvq���"��y5WP��9 �K�Oü���'���U�z"��lk����E^J��<��
��A�U��Q�Y�:�����&�t��}��Q ���b)N���G��&�铞E��� �+�>4�%�.���6�L&T1���������Ͳu㿋�TT6/<�$	�TK���y��X%�s���``Qo�n<�!������U�!Kp|�Ɖ�⌇=WeD�s�K!�J3b9���7�#�&����Fz��pI�I��]PK���<��QH�W�Sf��Ŀo����m7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3t��v'gn�]o��in�m��+�ވΦ�'�'�0�Xb�_�H�X�,\ަ�Itnh'yt�;U��֜��3�:ET֤vKzL͊�q����ϡ����pܜ!�I�lW���LWɆ&6�\]j}8o{:�֕ߝԀ�I�R���F��c��Z��}��	�d�bzP#�-������4Q��#��w21�X��|�C#/<���q��!�u�ǭ��k��?��}��7Q�� +@��牥��*[���Μ���a�M+|�����\��6fz5�WRj�.(Wx*q�\E��0�v�4�oK���-��%M�rs�i��UQA$��5�%]���a(􆿳����^���2jɸ�����5	���]���c�A�L'�������W��_�ړ8���/�}T���y~:���_EH��o��C!T*�q���U����?�!�`�(i3c��Et��q���U��;���)"����}���c��Et��q���U�ЂDa��(o��0��7c��Et��q���U��ꢤ�Og�ШT�7V��(�
t��Y�{'%s���䒼�W& s��Ѩg��U-�eE������(fx��V$�w�I�?g�f�;K�y��rk�gH��.��Fnt(L~΄gO�3��|��[��"�Q:�{�1hWw�d�pP;4��V�����q6�m��P��I��'�Po�Q�>�������IÙ=�HAmY�f��Ea�8Ss�LPo��p�(�oE��(��f��Q�m��'A>􏄃'�wZp�m~|��SpX�@>׼�\�v����ř�L�g?_��<'P��!jcCA�T�g�v����fQf��p�m~|����F}x�JHn��z�y���݈eG��{Ǧ%W& s���r7�����^���I���P4ǲ ���h9�5�܈zc��%��XP����c8?-+eN�Ȅ�4b�rS�b�8Z���'�e�����"�?;(��j67�Qs{ɯk�>p�m~|��7�q^�1�0M�/�s���'n�^0oy��\���W#�i'�6:	�<�&IMdK�Ch��T:���V�S�ff�݃зq8�Ј'���Xw�j�7��Po�Q�>°������R�wX��}�
�?�`<Y��sp4�r�@E�n`5�fK��0z�cULn�4Z_U���l�����"X��[��Q[R�7����n9읖w�x�z�f.�Э]�d�٣��c�A�L'�"��/f~�ƃ
ᾆ�x�T�\ ��i3�|)sՀ�T:���V����̵?oзq8�Ј'���Xw�j�7����;1�˚���ӯIJ ��`y����@����gG�������+N�f�+��Q]� _�rs�i�76b�*Ғ�ߨ�,R��g��U-�e,%�0g���l������*b��93��bj����Z鎬�������(������oD2��Я�R�wX��}�
�?�<��0n|�!h�b���t5a�l��0z�cULn�4Z_U���l����g��U-�e�j
��z�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��u�h����+Ed�J�5ٔ���)� ���2��5U`�������R�E�M��n��	�M�t%>^�ߡ�MQr��rY2r�b�@�|�S�Ժ��=�"��X��/c��!��q�=Ĉ���rl�$ho���<�n���p�n�����'�eEȆ���F1���\"��v��:�ߌ�JY�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���A����|������{,P�f�����t%>^�ߦ��|R%��<��0n|�!h�b���t-y|�$i�P�s+�¤]yFZ�%W�����8��'3��������h)C!nk��q-lC��ۺ_~W��8`ҧ��U�t����qE��6I&���#���i5�SKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hD}:��3��C����f�\� Iӥ�ѽ��L��[�1��4��}b2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �!-B=�6f�e9�R�[�̷��3hPo�Q�>°������R�wX�� �@��&}���$�K��=��Y�$���H&�4�1w<�?�ߨ�,R���"X��[�����D���G3҇
���2jɸx �M=�#����2jɸl
��������ӯIJ ��`y����T֣[\5g�1�9�U�WaU���|2s����ہ��!�#7ۏs|�L;Л�����V�M�$� %7䨹o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc<��H�M�6v�>%�fo C[�&x��`�ί�kG�X�`oò���?�~��-�Uٻ��
W⫃ ��5��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcu������MȆs��׾ŞWsuz'���Xw�j�7��AԢ�a\�T��}�%�`il��cf�p����b6vJ�pZ�*
T����}�r�KŸ���p�;����\uu�����r����!�`�(i3!�`�(i3Z鎬�������(����.��$�ʝ.�&J�!-B=�6f��c�t�{R��b�Bϱ�O�E�l`8x뛀���!���"��o_B�E�JQm��	�̷_��yC��S8�\�w�4�'�)�Բc��?!6)X���%A������D�ϲ]�6��2�S�i����T���!�`�(i3!�`�(i3!�`�(i3!�`�(i3��>��lJ���aٔ^?���S�T*��;1�˚�!��JlR����2jɸ\��)a�Pj �uw��o�Ķ
1'�F*�L��!�`�(i3!�`�(i3ouD�����rs�i� S�xSVe�W�6?��W��7(�bOpP�Fc�����k��$����导�?!6)X����*5���!�`�(i3!�`�(i3!�`�(i3!�`�(i36�&��=�'�)�Բck�A#�G=���%A������D�ϲ]�6��2Zb̶���~Lu��H�*b��93��/i�D���]�!��	Ǹ�y85��X��I�ՠ���aٔ^?��[+��.Ȉ�;1�˚�!��JlR�`<Y��sp(K�
�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3AԢ�a\����R�?�������|Pcsù�u�ȭ�>ѯN��S��I\�w[���!�`�(i3!�`�(i3!�`�(i3!�`�(i3-{�+2�p6ӆ�[W{b {��CWy)�+����$��r����!�`�(i3!�`�(i3Z鎬�������(����.��$��Z�d-�~E�`�_�y�1�����b��[� p!-B=�6f����k_!�`�(i3!�`�(i3!�`�(i3!�`�(i3X�o|3��b�Bϱ��!#��Rh�<Q�vn��l����I�/=k��%�W�%�K,�tc�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�2�~T����.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���߱QD�F�>u
���R ���q�l�:�r:���:�nl���~�?s5�b����c,�5<�'�ϖQֈE�^D��{�/�����v��M�0�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc]]� ?p�zw?��|��ՕH;u�o��_�Rv�䩲$���dS@Ɵ�o{y����i�q,?5q��C"�M��5�:��\���F�`yx�>�+X�[�G���K!�`�(i3!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}�D�wP�/�wۏ�:��"�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\��H����o�γ�ha��o���H�RtV�^xjzӝ�������iPo�Q�>��aIO-�����&G!�`�(i3p�n���/�i4?$|�ڗ�\���qhF�fp�Z��	�`D�\��v� H���;mQ��8���/���}Dq�f������!�`�(i3p�n���/�i4?$|�ڗ�\���x�o"jU�Z��	�`D�\��v� H���;mQ��8���/���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��C"�M�4��������L6�>P�2-i_m�;Y'�V!N�'�y�G